�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   Sexq0X   ChestPainTypeq1X	   RestingBPq2X   Cholesterolq3X	   FastingBSq4X
   RestingECGq5X   MaxHRq6etq7bX   n_features_in_q8KX
   n_outputs_q9KX   classes_q:h"h#K �q;h%�q<Rq=(KK�q>h)X   i8q?���q@RqA(KX   <qBNNNJ����J����K tqCb�C               qDtqEbX
   n_classes_qFKX   base_estimator_qGhX   estimators_qH]qI(h)�qJ}qK(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h8Kh9Kh:h"h#K �qLh%�qMRqN(KK�qOh)X   f8qP���qQRqR(KhBNNNJ����J����K tqSb�C              �?qTtqUbhFcnumpy.core.multiarray
scalar
qVhAC       qW�qXRqYX   max_features_qZKX   tree_q[csklearn.tree._tree
Tree
q\Kh"h#K �q]h%�q^Rq_(KK�q`hA�C       qatqbbK�qcRqd}qe(hKX
   node_countqfMWX   nodesqgh"h#K �qhh%�qiRqj(KMW�qkh)X   V56ql���qmRqn(Kh-N(X
   left_childqoX   right_childqpX   featureqqX	   thresholdqrX   impurityqsX   n_node_samplesqtX   weighted_n_node_samplesqutqv}qw(hoh)X   i8qx���qyRqz(KhBNNNJ����J����K tq{bK �q|hphzK�q}hqhzK�q~hrhRK�qhshRK �q�hthzK(�q�huhRK0�q�uK8KKtq�b�BK         ,                   @E@j8je3�?�           ��@       !                    �?P>�7���?L            @]@                          �Z@������?(             N@������������������������       �                     1@                          �Z@�lg����?            �E@������������������������       �                      @                           �?#z�i��?            �D@                          �_@�㙢�c�?             7@	                          �[@�IєX�?	             1@
                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     .@                            �?      �?             @������������������������       �                     �?                          @_@���Q��?             @������������������������       �                      @                          `b@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �c@X�<ݚ�?             2@                          �a@��S���?
             .@                            �?�q�q�?             "@������������������������       �                      @                          p`@և���X�?             @������������������������       �                     @������������������������       �                     @                          c@r�q��?             @                          �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @"       #                    �?0�)AU��?$            �L@������������������������       �                     G@$       +                   p`@�C��2(�?             &@%       *                    @z�G�z�?             @&       '                    �?      �?             @������������������������       �                      @(       )                    ]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @-       �                   �`@�ؗ���?�           H�@.       k                    �?��â�?�            �n@/       2                    �?H�g�}N�?v            �f@0       1                     �?��?^�k�?            �A@������������������������       �                     �?������������������������       �                     A@3       <                     �?
�n����?_            `b@4       9                   �p@      �?             0@5       6                    �?����X�?             @������������������������       �                     @7       8                   �^@      �?             @������������������������       �                      @������������������������       �                      @:       ;                   @_@�����H�?             "@������������������������       �                     �?������������������������       �                      @=       V                    �? ����?T            ``@>       ?                   �Q@���79��?=            @Y@������������������������       �                      @@       I                   0i@�C��2(�?<            �X@A       B                   `_@z�G�z�?             >@������������������������       �                     4@C       H                   �`@���Q��?             $@D       E                   �\@؇���X�?             @������������������������       �                     @F       G                    `@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @J       K                   @a@�nkK�?+            @Q@������������������������       �                     B@L       M                   @l@�C��2(�?            �@@������������������������       �                     &@N       S                    �?��2(&�?             6@O       R                   �a@�KM�]�?             3@P       Q                   @]@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             ,@T       U                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?W       Z                   �U@z�G�z�?             >@X       Y                    U@�q�q�?             @������������������������       �                     �?������������������������       �                      @[       j                    �?PN��T'�?             ;@\       e                   �`@����X�?             ,@]       d                    `@և���X�?             @^       c                   �^@���Q��?             @_       b                   �Z@�q�q�?             @`       a                   (q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @f       g                   �e@؇���X�?             @������������������������       �                     @h       i                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             *@l       �                    �?     ��?)             P@m       r                    �?�ՙ/�?             E@n       q                    ^@      �?              @o       p                     �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?s       �                    �?�t����?             A@t       �                    \@�������?             >@u       z                     �?��
ц��?	             *@v       y                   �u@�q�q�?             @w       x                   `X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @{       �                    Z@����X�?             @|       }                   @V@      �?             @������������������������       �                     �?~                          �X@�q�q�?             @������������������������       �                     �?�       �                   �j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�IєX�?             1@�       �                   �^@؇���X�?             @�       �                   @n@�q�q�?             @������������������������       �                     �?�       �                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�       �                   �_@      �?             @������������������������       �                     @������������������������       �                     �?�       �                     �?��2(&�?
             6@������������������������       �                     �?�       �                   @^@�����?	             5@������������������������       �                      @�       �                    �?8�Z$���?             *@������������������������       �                      @������������������������       �                     &@�       �                    �?��5��V�?�            0w@�       �                    �?Jܤm6�?;            �Y@�       �                     �?f.i��n�?            �F@�       �                   `a@������?	             1@�       �                   ``@�q�q�?             @������������������������       �                      @�       �                   �b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     &@�       �                   �Z@X�Cc�?             <@������������������������       �                      @�       �                   Pf@�	j*D�?             :@�       �                   �a@�}�+r��?             3@������������������������       �                     �?������������������������       �        
             2@������������������������       �                     @�       �                   �d@���y4F�?$            �L@�       �                   �l@$G$n��?            �B@������������������������       �                     *@�       �                   `d@�q�q�?             8@�       �                   �b@�㙢�c�?             7@�       �                    �?      �?              @�       �                   �b@����X�?             @�       �                    _@���Q��?             @������������������������       �                     �?�       �                   �q@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   �^@��S�ۿ?             .@�       �                   `]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?�       �                   �\@��Q��?             4@������������������������       �                     @�       �                     �?     ��?             0@������������������������       �                     @�       �                   Pe@�θ�?
             *@������������������������       �                     @�       �                    �?      �?              @�       �                   �h@      �?             @�       �                    d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    a@      �?             @������������������������       �                      @������������������������       �                      @�                          �?BO���V�?�            �p@�       �                    �?D��ٝ�?>            @Y@�       �                   �a@H�U?B�?2            �T@�       �                     �?4���C�?*            �P@�       �                   �Y@�eP*L��?             &@������������������������       �                      @�       �                   c@�q�q�?             "@�       �                   �p@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �\@r�q��?             @�       �                    k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   0c@���Q��?"            �K@�       �                   �b@V������?            �B@�       �                   0a@����"�?             =@�       �                    �?�	j*D�?             :@�       �                   �^@`�Q��?             9@�       �                   �[@�eP*L��?             &@������������������������       �                     �?�       �                   �a@      �?             $@�       �                   �o@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   `a@d}h���?             ,@������������������������       �                     @�       �                   �_@      �?              @������������������������       �                      @�       �                   �q@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   0d@b�2�tk�?             2@������������������������       �                     @�       �                   �`@��
ц��?             *@�       �                   �o@؇���X�?             @�       �                   �d@�q�q�?             @������������������������       �                     �?�       �                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �d@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   Xv@      �?             0@������������������������       �                     .@������������������������       �                     �?                         `@D�n�3�?             3@                        �]@�q�q�?             @                        �n@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @                          �?�	j*D�?             *@������������������������       �                      @                         a@���|���?             &@	      
                  ``@r�q��?             @������������������������       �                     �?������������������������       �                     @                        �b@���Q��?             @������������������������       �                     @������������������������       �                      @      4                  �`@r�q��?m             e@                        �a@�:�H:�?G            @[@                         @��s����?             5@                        Pa@z�G�z�?             4@������������������������       �                     &@                        �p@X�<ݚ�?             "@                         f@�q�q�?             @������������������������       �                     �?                        pa@z�G�z�?             @������������������������       �                      @                         �?�q�q�?             @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?       3                   @`���i��?9             V@!      *                   ]@Pq�����?7            @U@"      #                    �?@�0�!��?
             1@������������������������       �                      @$      )                   �?�q�q�?             "@%      &                  �l@      �?             @������������������������       �                      @'      (                  @[@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @+      2                   �? ��ʻ��?-             Q@,      -                  �p@@�E�x�?            �H@������������������������       �                     B@.      1                   d@$�q-�?             *@/      0                  �p@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     3@������������������������       �                     @5      B                  a@�k��(A�?&            �M@6      ?                   �?�eP*L��?             &@7      >                   �?�q�q�?             @8      9                  �b@���Q��?             @������������������������       �                     �?:      ;                    �?      �?             @������������������������       �                      @<      =                  Pi@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?@      A                  @q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?C      P                  �c@�q�q��?             H@D      M                   �?���Q��?             9@E      J                   �?�����?             3@F      G                   �?      �?
             0@������������������������       �                     $@H      I                  xp@�q�q�?             @������������������������       �                      @������������������������       �                     @K      L                  �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @N      O                  `c@�q�q�?             @������������������������       �                      @������������������������       �                     @Q      V                   b@�nkK�?             7@R      S                  `f@$�q-�?
             *@������������������������       �                     &@T      U                  ph@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KMWKK�q�hR�Bp       Ps@     �z@      1@      Y@      0@      F@              1@      0@      ;@       @              ,@      ;@      @      3@      �?      0@      �?      �?              �?      �?                      .@      @      @              �?      @       @       @              �?       @               @      �?              $@       @      @       @      @      @       @              @      @      @                      @      �?      @      �?       @               @      �?                      @      @              �?      L@              G@      �?      $@      �?      @      �?      @               @      �?      �?              �?      �?                      �?              @     @r@     Pt@     �J@      h@      8@     �c@      �?      A@      �?                      A@      7@      _@      @      $@      @       @      @               @       @       @                       @      �?       @      �?                       @      1@     �\@      &@     �V@       @              "@     �V@      @      8@              4@      @      @      @      �?      @              @      �?              �?      @                      @      @     �P@              B@      @      >@              &@      @      3@       @      1@       @      @       @                      @              ,@      �?       @               @      �?              @      8@       @      �?              �?       @              @      7@      @      $@      @      @      @       @      �?       @      �?      �?      �?                      �?              �?       @                       @      �?      @              @      �?      �?      �?                      �?              *@      =@     �A@      :@      0@       @      @      �?      @      �?                      @      �?              8@      $@      7@      @      @      @       @      @       @      �?              �?       @                      @      @       @       @       @      �?              �?       @              �?      �?      �?      �?                      �?      @              0@      �?      @      �?       @      �?      �?              �?      �?              �?      �?              @              $@              �?      @              @      �?              @      3@      �?               @      3@               @       @      &@       @                      &@     �m@     �`@     �M@     �E@      ,@      ?@      @      *@      @       @       @               @       @               @       @                      &@      $@      2@       @               @      2@      �?      2@      �?                      2@      @             �F@      (@      @@      @      *@              3@      @      3@      @      @      @      @       @      @       @      �?               @       @               @       @               @                      �?      ,@      �?      �?      �?      �?                      �?      *@                      �?      *@      @              @      *@      @      @              $@      @      @              @      @      @      �?      �?      �?      �?                      �?       @               @       @               @       @             �f@     @V@      D@     �N@      =@     �J@      <@      C@      @      @               @      @      @      �?       @      �?                       @      @      �?      �?      �?      �?                      �?      @              6@     �@@      &@      :@      &@      2@       @      2@       @      1@      @      @              �?      @      @      @      @      @                      @               @      @      &@              @      @      @               @      @      @              @      @                      �?      @                       @      &@      @      @              @      @      �?      @      �?       @              �?      �?      �?      �?                      �?              @      @      �?              �?      @              �?      .@              .@      �?              &@       @       @      @       @       @       @                       @               @      "@      @       @              @      @      @      �?              �?      @               @      @              @       @             �a@      <@     �X@      &@      1@      @      0@      @      &@              @      @       @      @      �?              �?      @               @      �?       @      �?      �?              �?      �?                      �?      @              �?             @T@      @     @T@      @      ,@      @       @              @      @      @      @       @              �?      @      �?                      @      @             �P@      �?      H@      �?      B@              (@      �?      @      �?              �?      @              @              3@                      @      E@      1@      @      @      @       @      @       @              �?      @      �?       @              �?      �?      �?                      �?      �?              �?      @              @      �?             �B@      &@      .@      $@      *@      @      (@      @      $@               @      @       @                      @      �?       @      �?                       @       @      @       @                      @      6@      �?      (@      �?      &@              �?      �?              �?      �?              $@        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfM=hgh"h#K �q�h%�q�Rq�(KM=�q�hn�BXE         *                   �^@4�5����?�           ��@                          `_@��hJ,�?V             a@       
                    a@��S�ۿ?%             N@       	                    �?�(\����?             D@                           �?Pa�	�?            �@@������������������������       �                     >@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                          �a@R���Q�?             4@������������������������       �                     @������������������������       �                     1@                          �`@���y4F�?1             S@                            �?�q�q�?             >@������������������������       �                      @                          0d@����X�?             <@                          c@�ՙ/�?             5@                          P`@������?             1@                           `@�r����?             .@                          �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             (@������������������������       �                      @������������������������       �                     @������������������������       �                     @                           �?�LQ�1	�?             G@������������������������       �                      @                          �\@��2(&�?             F@������������������������       �        
             *@        !                    ]@�n`���?             ?@������������������������       �                     @"       )                   �`@ �Cc}�?             <@#       $                    �?�S����?             3@������������������������       �                     @%       &                   �b@z�G�z�?	             .@������������������������       �                     $@'       (                   �c@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     "@+       �                   �`@4½D
��?s           ��@,       -                   �f@V^�b���?�            �l@������������������������       �        
             ,@.       }                    �?
Y�+ߧ�?�            �j@/       l                   �a@���_�?`             c@0       7                   �V@���U�?A            �Z@1       2                     �?�q�q�?             @������������������������       �                     �?3       6                    �?���Q��?             @4       5                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @8       9                    �?Ș����?=             Y@������������������������       �                     @@:       E                   �j@      �?,             Q@;       D                    �?��S���?	             .@<       =                   �[@���!pc�?             &@������������������������       �                     @>       ?                   �]@      �?              @������������������������       �                     �?@       A                    `@����X�?             @������������������������       �                      @B       C                   �h@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @F       G                    ]@�iʫ{�?#            �J@������������������������       �                     "@H       a                    �?�������?             F@I       ^                   �s@b�h�d.�?            �A@J       S                   �`@      �?             @@K       R                   �Z@�}�+r��?             3@L       M                   �o@؇���X�?             @������������������������       �                     @N       O                    _@      �?             @������������������������       �                      @P       Q                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@T       U                     �?�θ�?	             *@������������������������       �                     @V       W                   0a@�q�q�?             "@������������������������       �                     �?X       ]                    �?      �?              @Y       Z                   �k@؇���X�?             @������������������������       �                     @[       \                    ]@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?_       `                     �?�q�q�?             @������������������������       �                      @������������������������       �                     �?b       k                    �?�q�q�?             "@c       d                   Pk@և���X�?             @������������������������       �                     �?e       j                   @^@�q�q�?             @f       g                     �?�q�q�?             @������������������������       �                     �?h       i                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @m       r                     �?dP-���?            �G@n       o                   �^@      �?             @������������������������       �                     �?p       q                   Xs@�q�q�?             @������������������������       �                      @������������������������       �                     �?s       t                   �[@ �#�Ѵ�?            �E@������������������������       �                     6@u       v                   �c@�����?             5@������������������������       �        	             ,@w       x                    ]@����X�?             @������������������������       �                     �?y       |                   �q@r�q��?             @z       {                   �m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @~       �                   �`@      �?,             O@       �                   �Z@���y4F�?             3@�       �                   @_@�q�q�?             @������������������������       �                     @�       �                   �X@�q�q�?             @������������������������       �                     �?�       �                     �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             *@�       �                    �?�lg����?            �E@�       �                    k@8�A�0��?             6@������������������������       �                     "@�       �                   �o@�	j*D�?             *@�       �                   `m@      �?              @�       �                    �?z�G�z�?             @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?؇���X�?             5@������������������������       �                     �?�       �                   8r@ףp=
�?             4@������������������������       �        
             0@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?��5��?�            w@�       �                    �?fC�K�q�?J             `@�       �                   �p@�����?             C@�       �                   �j@      �?             2@������������������������       �                     @�       �                   �c@�	j*D�?             *@�       �                   �a@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �`@R���Q�?	             4@������������������������       �                     "@�       �                   xu@���!pc�?             &@������������������������       �                     @�       �                   y@      �?             @������������������������       �                     @������������������������       �                     @�       �                     �?fK!���?6            �V@�       �                    �?���Q��?
             4@�       �                    c@�t����?             1@�       �                    b@����X�?             @�       �                   �l@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     $@������������������������       �                     @�       �                   �b@X3_��?,            �Q@�       �                   �a@�G\�c�?(            @P@�       �                    g@V{q֛w�?&             O@�       �                   �e@�C��2(�?             &@������������������������       �                     @�       �                   `c@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?!            �I@�       �                   �b@�I� �?             G@�       �                   @b@\X��t�?             7@�       �                    �?8�A�0��?             6@�       �                   �o@�z�G��?             $@�       �                    _@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    a@      �?             (@�       �                   @^@؇���X�?             @�       �                   �n@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   @c@��<b���?             7@������������������������       �                     @�       �                   �t@     ��?
             0@�       �                   pd@d}h���?	             ,@�       �                   �c@      �?             @������������������������       �                     �?�       �                   �]@���Q��?             @������������������������       �                     �?�       �                   �k@      �?             @������������������������       �                      @�       �                   d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   `a@���Q��?             @������������������������       �                     �?�       �                   �]@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �b@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                     �?�Q��k�?�             n@�       �                   �c@ Df@��?/            �T@�       �                   0h@@4և���?             <@������������������������       �                      @������������������������       �                     :@������������������������       �                    �K@�       �                   pi@�xV�w�?d            �c@�       �                   �g@�}�+r��?             C@�       �                    �?�����?             5@������������������������       �                     @�       �                   `^@      �?
             0@������������������������       �                     �?�       �                   a@��S�ۿ?	             .@�       �                    �?r�q��?             @�       �                   @e@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     1@�       :                   �?�t����?O            �]@�       +                  e@����x�?I            @[@�       (                   �?�û��|�?/            @Q@�                          �?      �?+             P@�                         @o@�����?             3@                          @     ��?
             0@                        �\@      �?             (@                        `m@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @      	                  `a@���Q��?            �F@������������������������       �                     @
      '                   t@�\��N��?             C@      &                  8r@X�<ݚ�?             B@                        �`@��.k���?             A@                        �a@��H�}�?             9@������������������������       �                     @                        �l@���!pc�?             6@������������������������       �                     @                        �l@ҳ�wY;�?             1@������������������������       �                      @                         q@������?
             .@                        �^@���|���?             &@                        �b@և���X�?             @                        0m@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        �o@      �?             @                        �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @       %                  �d@�<ݚ�?             "@!      $                   �?      �?              @"      #                   b@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @)      *                  @_@���Q��?             @������������������������       �                      @������������������������       �                     @,      9                   f@z�G�z�?             D@-      2                   m@������?            �B@.      /                   �?և���X�?             @������������������������       �                     @0      1                  �`@      �?             @������������������������       �                     @������������������������       �                     �?3      4                   �?(;L]n�?             >@������������������������       �                     5@5      8                   f@�����H�?             "@6      7                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @;      <                  �k@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@q�tq�bh�h"h#K �q�h%�q�Rq�(KM=KK�q�hR�B�       �t@     y@      4@      ]@      @      L@      �?     �C@      �?      @@              >@      �?       @      �?                       @              @      @      1@      @                      1@      0@      N@      $@      4@       @               @      4@       @      *@      @      *@       @      *@       @      �?              �?       @                      (@       @              @                      @      @      D@               @      @      C@              *@      @      9@      @              @      9@      @      0@              @      @      (@              $@      @       @      @                       @              "@     �s@     �q@      L@     �e@              ,@      L@     �c@      9@      `@      5@     @U@      @       @      �?              @       @      �?       @               @      �?               @              1@     �T@              @@      1@     �I@       @      @       @      @      @              @      @              �?      @       @       @              @       @      @                       @              @      "@      F@              "@      "@     �A@      @      =@      @      <@      �?      2@      �?      @              @      �?      @               @      �?      �?      �?                      �?              (@      @      $@              @      @      @      �?               @      @      �?      @              @      �?      @      �?                      @      �?               @      �?       @                      �?      @      @      @      @      �?               @      @       @      �?      �?              �?      �?      �?                      �?              @               @      @     �E@       @       @              �?       @      �?       @                      �?       @     �D@              6@       @      3@              ,@       @      @      �?              �?      @      �?       @               @      �?                      @      ?@      ?@      .@      @       @      @              @       @      �?      �?              �?      �?              �?      �?              *@              0@      ;@      *@      "@      "@              @      "@      @      @      �?      @      �?      �?              �?      �?                      @      @                      @      @      2@      �?               @      2@              0@       @       @       @                       @     p@      \@      L@     @R@      (@      :@      "@      "@              @      "@      @      �?      @      �?                      @       @              @      1@              "@      @       @              @      @      @      @                      @      F@     �G@      (@       @      (@      @       @      @       @       @       @                       @              @      $@                      @      @@     �C@      ;@      C@      ;@     �A@      $@      �?      @              @      �?      @                      �?      1@      A@      .@      ?@      $@      *@      "@      *@      @      @      @      �?      @                      �?              @      @      @      @      �?      @      �?      @                      �?      �?                      @      �?              @      2@              @      @      &@      @      &@      @      @      �?               @      @      �?              �?      @               @      �?      �?      �?                      �?               @       @               @      @      �?              �?      @      �?                      @              @      @      �?      @                      �?      i@     �C@     @T@       @      :@       @               @      :@             �K@              ^@     �B@      B@       @      3@       @      @              ,@       @              �?      ,@      �?      @      �?       @      �?              �?       @              @              "@              1@              U@     �A@     �R@      A@      E@      ;@      D@      8@      *@      @      *@      @      "@      @      �?      @              @      �?               @              @                      @      ;@      2@      @              4@      2@      4@      0@      2@      0@      0@      "@              @      0@      @      @              &@      @               @      &@      @      @      @      @      @       @      �?       @                      �?      �?      @      �?      �?              �?      �?                       @      @              @               @      @      �?      @      �?      @      �?                      @              @      �?               @                       @       @      @       @                      @     �@@      @     �@@      @      @      @      @              �?      @              @      �?              =@      �?      5@               @      �?      �?      �?              �?      �?              @                      @      "@      �?              �?      "@        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfM=hgh"h#K �q�h%�q�Rq�(KM=�q�hn�BXE                              _@p�Vv���?�           ��@                          `\@D��*�4�?^            @a@������������������������       �        #             K@                           �?���H��?;             U@                           �?(;L]n�?)             N@                           �?�t����?             1@������������������������       �                     @       	                    `@z�G�z�?             $@������������������������       �                     �?
                          �b@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                    �E@                           @�q�q�?             8@                           �?D�n�3�?             3@                            �?�eP*L��?	             &@������������������������       �                     �?                          �]@      �?             $@������������������������       �                     @                           `@r�q��?             @������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?      �?              @                          �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          p`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @!       R                     �?n��mb��?�           ��@"       Q                   Pe@�g+�v�?S             a@#       >                    �?�"'`�]�?E            @\@$       -                   �_@<|ۤ$�?            �K@%       ,                    �?���!pc�?
             6@&       )                   �p@�q�q�?	             2@'       (                   �`@d}h���?             ,@������������������������       �                     &@������������������������       �                     @*       +                    `@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @.       ;                   �u@�'�`d�?            �@@/       :                   �e@r�q��?             >@0       5                   �a@\-��p�?             =@1       2                   @]@�q�q�?             "@������������������������       �                      @3       4                   @b@؇���X�?             @������������������������       �                     @������������������������       �                     �?6       9                   Pp@P���Q�?             4@7       8                   @o@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?<       =                   0c@�q�q�?             @������������������������       �                     �?������������������������       �                      @?       B                    [@�8���?&             M@@       A                   �m@�q�q�?             @������������������������       �                      @������������������������       �                     �?C       D                    �?h㱪��?$            �K@������������������������       �                     =@E       F                   @a@$�q-�?             :@������������������������       �                     $@G       P                    �?      �?	             0@H       O                    @�r����?             .@I       L                   �a@"pc�
�?             &@J       K                   Pn@�q�q�?             @������������������������       �                      @������������������������       �                     �?M       N                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     7@S                          xp@b �>��?.           �|@T       �                   �`@���f��?�            �t@U       V                   `Z@ �]^m>�?{             g@������������������������       �                     @W       �                    �?�K��?w            @f@X       �                   ``@��=A��?8             S@Y       �                    �?ҳ�wY;�?4             Q@Z       y                   d@l��
I��?+             K@[       l                   �\@��|�5��?&            �G@\       _                    �?�n_Y�K�?             *@]       ^                   @k@      �?             @������������������������       �                      @������������������������       �                      @`       k                   �o@�q�q�?	             "@a       j                    �?և���X�?             @b       i                   �n@�q�q�?             @c       h                   @a@z�G�z�?             @d       e                   `_@�q�q�?             @������������������������       �                     �?f       g                   �k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @m       t                    g@@�0�!��?             A@n       o                   �`@�n_Y�K�?             *@������������������������       �                     @p       s                   @_@����X�?             @q       r                   �a@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @u       v                   �_@���N8�?             5@������������������������       �        	             $@w       x                   Hp@�C��2(�?	             &@������������������������       �                     $@������������������������       �                     �?z       {                   �i@����X�?             @������������������������       �                     �?|       }                   �d@r�q��?             @������������������������       �                     @~                           k@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �_@և���X�?	             ,@�       �                   �_@����X�?             @������������������������       �                      @�       �                   �n@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    `@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                   `a@��x_F-�??            �Y@�       �                   �Z@ܷ��?��?             =@�       �                   `V@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �? �q�q�?             8@������������������������       �                     @�       �                    `@�X�<ݺ?	             2@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                   �l@x�� ���?/            @R@�       �                   `d@�LQ�1	�?             G@�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @�ʈD��?            �E@�       �                    �?@4և���?             E@������������������������       �                     ;@�       �                   ``@z�G�z�?
             .@�       �                   `j@؇���X�?	             ,@������������������������       �                     "@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   `m@�5��?             ;@�       �                   pc@؇���X�?             @�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?      �?             4@�       �                   �o@������?             1@�       �                    c@ףp=
�?             $@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �_@և���X�?             @�       �                   �^@���Q��?             @�       �                   �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �b@H�+��<�?`            �b@�       �                    �?\������?E            @Z@�       �                   �h@���-T��?*             O@�       �                   �^@���Q��?
             .@������������������������       �                     "@������������������������       �                     @�       �                    �?=QcG��?             �G@�       �                   �k@����X�?             @������������������������       �                     @�       �                   `c@      �?             @������������������������       �                     �?�       �                   `_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�(\����?             D@�       �                   �b@(;L]n�?             >@������������������������       �                     0@�       �                   �`@@4և���?	             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �        
             $@�       �                   @j@v ��?            �E@�       �                    [@�q�q�?	             .@������������������������       �                     @�       �                   `c@r�q��?             (@�       �                    �?����X�?             @������������������������       �                     @�       �                   b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?X�Cc�?             <@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     @�       �                   pb@      �?             4@�       �                   o@�8��8��?             (@������������������������       �                      @�       �                   �a@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   m@      �?              @�       �                    k@z�G�z�?             @�       �                    X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   `f@�GN�z�?             F@�       �                   `d@$G$n��?            �B@�       �                   �j@�t����?
             1@�       �                   c@�eP*L��?             &@������������������������       �                     @�       �                   �f@      �?              @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     4@�       �                   �l@����X�?             @������������������������       �                     @������������������������       �                      @                        Hq@�U���?S            �_@      	                  �`@��]�T��?            �D@                         �?�}�+r��?             3@                        8q@��S�ۿ?             .@������������������������       �        	             *@                        �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @
                        0c@���|���?             6@                         �?X�<ݚ�?             "@                         �?      �?              @                        �`@z�G�z�?             @                        Pb@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?                          @�θ�?             *@                        �p@r�q��?             (@������������������������       �                     @                        �p@      �?              @������������������������       �                     �?                        �d@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?      2                  �s@&^�)b�?7            �U@      -                  `e@      �?(             P@                         @a@�U�:��?#            �M@������������������������       �                     7@!      ,                  Hr@4?,R��?             B@"      '                   �?���N8�?             5@#      &                  �q@ףp=
�?             $@$      %                  �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @(      )                   �?���|���?             &@������������������������       �                      @*      +                  pb@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     .@.      1                   �?���Q��?             @/      0                  �q@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?3      <                  c@���|���?             6@4      9                   �?��.k���?             1@5      6                   �?z�G�z�?             $@������������������������       �                     @7      8                  v@�q�q�?             @������������������������       �                     �?������������������������       �                      @:      ;                  @[@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @q�tq�bh�h"h#K �q�h%�q�Rq�(KM=KK�q�hR�B�       @t@     �y@      $@      `@              K@      $@     �R@       @      M@       @      .@              @       @       @      �?              �?       @               @      �?                     �E@       @      0@       @      &@      @      @      �?              @      @      @              �?      @              @      �?      �?      �?                      �?       @      @      �?       @      �?                       @      �?      @      �?                      @              @     �s@     �q@     @Y@     �A@     �S@     �A@      7@      @@      0@      @      (@      @      &@      @      &@                      @      �?      @      �?                      @      @              @      :@      @      9@      @      9@      @      @       @              �?      @              @      �?              �?      3@      �?      @              @      �?                      *@      �?               @      �?              �?       @             �K@      @       @      �?       @                      �?     �J@       @      =@              8@       @      $@              ,@       @      *@       @      "@       @       @      �?       @                      �?      @      �?      @                      �?      @              �?              7@             �j@     �n@     �f@     �b@     �]@     @P@      @             @\@     @P@      ?@     �F@      8@      F@      0@      C@      &@      B@      @       @       @       @       @                       @      @      @      @      @       @      @      �?      @      �?       @              �?      �?      �?      �?                      �?               @      �?              �?                       @      @      <@      @       @              @      @       @      @       @      @                       @       @              �?      4@              $@      �?      $@              $@      �?              @       @              �?      @      �?      @               @      �?              �?       @               @      @      @       @       @              @       @      @                       @      @      @      @                      @      @      �?              �?      @             �T@      4@      :@      @      @       @      @                       @      7@      �?      @              1@      �?      @      �?      @                      �?      $@              L@      1@      D@      @      �?       @      �?                       @     �C@      @     �C@      @      ;@              (@      @      (@       @      "@              @       @      @                       @              �?              �?      0@      &@      �?      @      �?       @      �?                       @              @      .@      @      *@      @      "@      �?       @      �?      �?              �?      �?              �?      �?              @              @      @       @      @       @      �?              �?       @                       @       @               @      �?              �?       @             �O@     �U@      =@      S@      "@     �J@      @      "@              "@      @              @      F@       @      @              @       @       @              �?       @      �?              �?       @              �?     �C@      �?      =@              0@      �?      *@              *@      �?                      $@      4@      7@      $@      @              @      $@       @      @       @      @              �?       @      �?                       @      @              $@      2@      @      @      @                      @      @      .@      �?      &@               @      �?      @      �?                      @      @      @      �?      @      �?      �?              �?      �?                      @      @              A@      $@      @@      @      (@      @      @      @      @              @      @      @      �?              �?      @                      @      @              4@               @      @              @       @              ?@      X@      .@      :@      �?      2@      �?      ,@              *@      �?      �?      �?                      �?              @      ,@       @      @      @      @      @      �?      @      �?       @      �?                       @               @      @                      �?      $@      @      $@       @      @              @       @              �?      @      �?      @                      �?              �?      0@     �Q@       @      L@      @      K@              7@      @      ?@      @      0@      �?      "@      �?      �?              �?      �?                       @      @      @               @      @      @      @                      @              .@      @       @      @      �?              �?      @                      �?       @      ,@       @      "@       @       @              @       @      �?              �?       @              @      �?              �?      @                      @q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       qՆq�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}q�(hKhfM+hgh"h#K �q�h%�q�Rq�(KM+�q�hn�BhA                            �?U�ք�?�           ��@       3                   �c@^��I��?u           ��@                            �?ڤ���?4            @T@                          �Z@$gv&��?&            �M@������������������������       �                     @                            �?�T`�[k�?#            �J@������������������������       �                     @                           `@j�q����?              I@	                           I@��p\�?            �D@
                          �]@��a�n`�?             ?@                           �?     ��?             0@������������������������       �                      @                           �?d}h���?
             ,@                          p`@      �?              @                           �?�q�q�?             @                          �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          @\@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     .@������������������������       �                     $@                           b@�q�q�?             "@                          @E@؇���X�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @!       2                   `Q@���|���?             6@"       1                   @e@�q�q�?             5@#       $                     �?�d�����?             3@������������������������       �                     �?%       (                   �_@�E��ӭ�?             2@&       '                   �[@      �?             @������������������������       �                     �?������������������������       �                     @)       .                    �?؇���X�?             ,@*       +                   `b@�C��2(�?             &@������������������������       �                     @,       -                   �c@      �?             @������������������������       �                     �?������������������������       �                     @/       0                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?4       �                    �?��S�[�?A            ~@5       �                   �e@V������?�            �k@6       m                   �`@�d�����?�             j@7       Z                    �?      �?J             \@8       S                    `@�)V���?;            @V@9       F                   pj@F.< ?�?.            �P@:       ;                     �?p�ݯ��?             3@������������������������       �                     �?<       =                   @_@�q�q�?             2@������������������������       �                     @>       E                   �h@      �?
             (@?       @                   �\@      �?              @������������������������       �                     @A       D                   �a@���Q��?             @B       C                   pg@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @G       R                   �a@��E�B��?            �G@H       Q                   �a@     ��?             @@I       J                   `p@ܷ��?��?             =@������������������������       �                     5@K       P                   �`@      �?              @L       M                     �?����X�?             @������������������������       �                     �?N       O                   �p@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        	             .@T       U                     �?
;&����?             7@������������������������       �                     $@V       W                    �?8�Z$���?             *@������������������������       �                     @X       Y                   �j@����X�?             @������������������������       �                      @������������������������       �                     @[       ^                     �?��+7��?             7@\       ]                   @_@      �?             @������������������������       �                     @������������������������       �                     �?_       d                   �[@�d�����?             3@`       a                   @_@      �?              @������������������������       �                     �?b       c                   �n@؇���X�?             @������������������������       �                     @������������������������       �                     �?e       j                   �^@���|���?             &@f       g                    ]@      �?             @������������������������       �                      @h       i                   �\@      �?             @������������������������       �                     @������������������������       �                     �?k       l                   �k@z�G�z�?             @������������������������       �                     �?������������������������       �                     @n       �                   pn@�*v��?@            @X@o       �                    �?�����?!            �H@p       �                   `l@���?            �D@q       x                   �h@6YE�t�?            �@@r       s                     �?�q�q�?             "@������������������������       �                     �?t       u                   @a@      �?              @������������������������       �                      @v       w                   �`@r�q��?             @������������������������       �                     @������������������������       �                     �?y       z                   �Y@�8��8��?             8@������������������������       �                     �?{       �                   �j@�nkK�?             7@|       }                   �b@�����H�?             "@������������������������       �                     @~                          �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@�       �                     �?      �?              @������������������������       �                     �?�       �                   �a@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                   pd@      �?             H@�       �                    �?����?�?            �F@������������������������       �                    �A@�       �                   �p@ףp=
�?             $@������������������������       �                     @�       �                   �]@z�G�z�?             @������������������������       �                     @�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   pe@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �f@8�Z$���?             *@�       �                     �?�q�q�?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?�       �                   l@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   @\@<�I<���?�             p@�       �                    g@D�n�3�?             3@�       �                     �?ҳ�wY;�?             1@�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�n_Y�K�?	             *@�       �                   @\@      �?             $@������������������������       �                     �?�       �                    �?X�<ݚ�?             "@�       �                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �X@      �?             @������������������������       �                     �?�       �                    �?���Q��?             @������������������������       �                      @�       �                   @e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                     �?R7�#�z�?�            �m@�       �                   `c@�(\����?6             T@�       �                   �q@�"w����?3             S@������������������������       �        (            �O@�       �                   0r@$�q-�?             *@������������������������       �                     �?������������������������       �        
             (@�       �                   @e@      �?             @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   pl@�N����?k            �c@�       �                   ``@l��\��?,             Q@�       �                   �_@�(\����?             D@������������������������       �                     <@�       �                    �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?�       �                   Pi@�>4և��?             <@�       �                   �`@P���Q�?             4@�       �                   `e@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             .@�       �                   Pa@      �?              @������������������������       �                     @�       �                   �k@z�G�z�?             @������������������������       �                      @�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   Pm@��|�	��??            �V@�       �                    @�����?
             3@�       �                   �c@և���X�?             ,@�       �                    _@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �l@����X�?             @������������������������       �                     @�       �                    b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�                         �d@      �?5             R@�       �                   `]@H�V�e��?3             Q@�       �                   `\@      �?              @�       �                   �Z@�q�q�?             @������������������������       �                     �?�       �                    @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                   �c@r�q��?.             N@�       �                   pa@�z�G��?             >@�       �                    @@4և���?             ,@������������������������       �        
             *@������������������������       �                     �?�       �                    �?      �?             0@�       �                    b@      �?              @������������������������       �                      @�       �                    �?�q�q�?             @�       �                   �q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �`@      �?              @�       �                    @      �?             @�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�                           �?(;L]n�?             >@�       �                   �d@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     7@������������������������       �                     @                         �?H~4o]�?j            �e@                        �p@Hn�.P��?J             _@������������������������       �        =            �Y@                        �_@����X�?             5@                        c@      �?             (@                         �?�q�q�?             "@	      
                  �S@���Q��?             @������������������������       �                     �?                        �Z@      �?             @������������������������       �                     �?                        �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     "@      &                  �b@Tt�ó��?             �H@      %                  pr@�'�`d�?            �@@                        �`@�חF�P�?             ?@                         �?P���Q�?             4@                        �Y@      �?              @                        �W@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     (@      $                  0o@���|���?	             &@                         �?և���X�?             @������������������������       �                     �?       !                   �?      �?             @������������������������       �                      @"      #                  `^@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @'      (                  �e@      �?
             0@������������������������       �                     &@)      *                  �p@z�G�z�?             @������������������������       �                     @������������������������       �                     �?q�tq�bh�h"h#K �q�h%�q�Rq�(KM+KK�q�hR�B�        t@     �y@     `r@     �p@      4@     �N@      (@     �G@              @      (@     �D@      @              "@     �D@      @      C@      @      <@      @      *@               @      @      &@      �?      @      �?       @      �?      �?              �?      �?                      �?              @       @      @              @       @                      .@              $@      @      @      @      �?      �?      �?              �?      �?              @                       @       @      ,@      @      ,@      @      ,@              �?      @      *@      @      �?              �?      @               @      (@      �?      $@              @      �?      @      �?                      @      �?       @      �?                       @       @              �?              q@     �i@     �P@     �c@     �K@     @c@      E@     �Q@      9@      P@      *@     �J@      @      (@      �?              @      (@              @      @      @       @      @              @       @      @       @      �?       @                      �?               @      @              @     �D@      @      :@      @      :@              5@      @      @       @      @      �?              �?      @      �?                      @      �?              @                      .@      (@      &@      $@               @      &@              @       @      @       @                      @      1@      @      @      �?      @                      �?      ,@      @      @      �?      �?              @      �?      @                      �?      @      @      @      @               @      @      �?      @                      �?      @      �?              �?      @              *@      U@      $@     �C@      $@      ?@      @      <@      @      @              �?      @      @       @              �?      @              @      �?               @      6@      �?              �?      6@      �?       @              @      �?      �?      �?                      �?              ,@      @      @              �?      @       @      @                       @               @      @     �F@      �?      F@             �A@      �?      "@              @      �?      @              @      �?      �?      �?                      �?       @      �?       @                      �?      &@       @      @       @       @               @       @              �?       @      �?              �?       @              @              j@      I@       @      &@      @      &@      �?      @              @      �?              @       @      @      @      �?              @      @      �?       @      �?                       @      @      @              �?      @       @       @              �?       @               @      �?                      @       @              i@     �C@     �S@       @     �R@      �?     �O@              (@      �?              �?      (@              @      �?      �?      �?      �?                      �?       @             �^@     �B@      O@      @     �C@      �?      <@              &@      �?      &@                      �?      7@      @      3@      �?      @      �?              �?      @              .@              @      @              @      @      �?       @               @      �?              �?       @              N@      ?@      @      *@      @       @      @      @      @                      @       @      @              @       @       @               @       @                      @      K@      2@      K@      ,@      @      @      @       @      �?              @       @      @                       @               @      I@      $@      5@      "@      *@      �?      *@                      �?       @       @      @       @       @              @       @      @      �?      @                      �?              �?       @      @       @       @       @      �?              �?       @                      �?              @      =@      �?      @      �?              �?      @              7@                      @      <@      b@      @     �]@             �Y@      @      .@      @      @      @      @      @       @      �?               @       @              �?       @      �?              �?       @                      @      @                      "@      6@      ;@      @      :@      @      :@      �?      3@      �?      @      �?      �?              �?      �?                      @              (@      @      @      @      @      �?              @      @       @              �?      @              @      �?                      @       @              .@      �?      &@              @      �?      @                      �?q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h8Kh9Kh:h"h#K �q�h%�q�Rq�(KK�q�hR�C              �?q�tq�bhFhVhAC       q��q�Rq�hZKh[h\Kh"h#K �q�h%�q�Rq�(KK�q�hA�C       q�tq�bK�q�Rq�}r   (hKhfMOhgh"h#K �r  h%�r  Rr  (KMO�r  hn�BHI         �                   �`@4�5����?�           ��@       o                    �?��#e���?�            �t@       >                    �?>����|�?�            �m@       #                    �?�A��c�?j            `e@                           `_@hdpZ�L�?K            @\@                          �[@��<D�m�??            �X@                            �?�q��/��?             G@       	                   �X@���Q��?             @������������������������       �                     �?
                          �p@      �?             @������������������������       �                     @������������������������       �                     �?                          �a@��p\�?            �D@                          `[@ȵHPS!�?             :@                          �o@P���Q�?             4@������������������������       �                     &@                           �?�����H�?             "@������������������������       �                     @                          �p@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                          �j@�q�q�?             @������������������������       �                     @                          �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             .@                           _@ pƵHP�?!             J@������������������������       �                     F@                            �?      �?              @������������������������       �                     �?������������������������       �                     @!       "                   j@���Q��?             .@������������������������       �                     @������������������������       �                     "@$       1                   �`@����"�?             M@%       (                     �?X�<ݚ�?             ;@&       '                   pj@���Q��?             @������������������������       �                      @������������������������       �                     @)       0                   �q@�eP*L��?             6@*       /                    `@p�ݯ��?
             3@+       .                   �Y@�t����?	             1@,       -                   `Z@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@������������������������       �                      @������������������������       �                     @2       9                   �e@��a�n`�?             ?@3       8                   @`@�LQ�1	�?             7@4       7                    S@�C��2(�?             6@5       6                   @b@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@������������������������       �                     �?:       ;                     �?      �?              @������������������������       �                     @<       =                   �q@z�G�z�?             @������������������������       �                     @������������������������       �                     �??       n                   �_@����e��?0            �P@@       m                    g@|��?���?*             K@A       f                    �?�q�����?)             I@B       E                   �Z@��Zy�?             �C@C       D                   �Z@z�G�z�?             @������������������������       �                     �?������������������������       �                     @F       K                     �?h+�v:�?             A@G       J                   @e@�<ݚ�?             "@H       I                   `Z@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?L       W                   c@� �	��?             9@M       R                    �?�q�q�?             "@N       O                   Pb@      �?             @������������������������       �                     �?P       Q                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?S       T                   @\@z�G�z�?             @������������������������       �                     @U       V                   `^@      �?              @������������������������       �                     �?������������������������       �                     �?X       [                   �X@     ��?             0@Y       Z                   `V@      �?             @������������������������       �                     �?������������������������       �                     @\       a                   @[@r�q��?             (@]       ^                    a@�q�q�?             @������������������������       �                     �?_       `                   @d@      �?              @������������������������       �                     �?������������������������       �                     �?b       c                   �]@�����H�?             "@������������������������       �                     @d       e                    �?      �?             @������������������������       �                     �?������������������������       �                     @g       l                    �?"pc�
�?	             &@h       i                   �`@�q�q�?             @������������������������       �                     �?j       k                    c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     (@p       �                   Pz@     ��?E             X@q       x                     �?heu+��?D            �W@r       s                   �Y@      �?              @������������������������       �                     @t       w                   `^@z�G�z�?             @u       v                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @y       |                    �?��+��<�?=            �U@z       {                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?}       ~                   pa@F|/ߨ�?8            @T@������������������������       �        !             G@       �                    �? >�֕�?            �A@�       �                   �a@8�Z$���?
             *@�       �                   @a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �\@�C��2(�?             &@�       �                    [@      �?             @������������������������       �                      @�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     6@������������������������       �                      @�                         d@>@��?           y@�       �                   @E@n�QJ���?�            `o@�       �                    �?\-��p�?             =@�       �                    _@���7�?             6@�       �                    �?      �?              @�       �                     �?r�q��?             @������������������������       �                     @�       �                   `]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@�       �                   pb@և���X�?             @�       �                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �n@` .�(�?�            �k@�       �                   �`@J��	�y�?S            @_@�       �                    �?0,Tg��?6             U@�       �                    �?     ��?,             P@�       �                   �b@�G�z��?             4@�       �                    a@d}h���?
             ,@������������������������       �                     �?�       �                     �?8�Z$���?	             *@������������������������       �                     @�       �                   �m@z�G�z�?             $@�       �                   �j@�����H�?             "@������������������������       �                     @�       �                   `]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?t��ճC�?             F@������������������������       �                     0@�       �                   `b@ �Cc}�?             <@������������������������       �        	             *@�       �                   �l@z�G�z�?	             .@������������������������       �                     (@������������������������       �                     @�       �                    �?      �?
             4@�       �                   �j@      �?             0@������������������������       �                     @�       �                    �?�q�q�?             "@�       �                    \@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   Pf@v�2t5�?            �D@�       �                    �?      �?              @�       �                   0a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�'�=z��?            �@@�       �                   pj@�f7�z�?             =@�       �                   �h@      �?              @������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                      @�       �                   �i@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    a@����X�?             5@�       �                   c@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �k@�r����?             .@������������������������       �                     @�       �                    �?"pc�
�?	             &@�       �                   �a@ףp=
�?             $@������������������������       �                     @�       �                   �b@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�{<����?=            @X@�       �                    �?r�qG�?              H@�       �                    f@�7����?            �G@�       �                    �?��Hg���?            �F@�       �                    b@�GN�z�?             F@�       �                   �`@�q�q�?             5@�       �                   �o@      �?             ,@������������������������       �                     @�       �                   xp@���|���?             &@������������������������       �                     @�       �                   8s@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    q@�LQ�1	�?             7@������������������������       �                     $@�       �                   Pq@�θ�?
             *@������������������������       �                     �?�       �                     �?r�q��?	             (@�       �                   pc@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �p@`�(c�?            �H@�       �                   @o@z�G�z�?             .@������������������������       �                     �?�       �                   �b@؇���X�?             ,@������������������������       �                     $@�       �                    �?      �?             @�       �                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?                         �c@H�V�e��?             A@                        �b@HP�s��?             9@                        `c@؇���X�?
             ,@������������������������       �                     (@������������������������       �                      @������������������������       �                     &@                        |@X�<ݚ�?             "@                        �\@����X�?             @������������������������       �                     �?	      
                  �c@r�q��?             @������������������������       �                     @                        �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @      F                   �?H.�!���?b            �b@      E                  @g@�+$�jP�?W            �`@      &                   �?�{�@�N�?V            �`@                        �i@��>4և�?             <@������������������������       �                     @                        �p@`�Q��?             9@                        �k@�8��8��?
             (@������������������������       �                     @                        �b@r�q��?             @������������������������       �                     @������������������������       �                     �?                          �?��
ц��?             *@������������������������       �                     @                         ^@���Q��?             $@������������������������       �                     @      %                  0f@�q�q�?             @                         �`@z�G�z�?             @������������������������       �                      @!      "                   �?�q�q�?             @������������������������       �                     �?#      $                  pe@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?'      ,                   �?(N:!���?B            @Z@(      +                  m@(;L]n�?#             N@)      *                  `l@$�q-�?             :@������������������������       �                     8@������������������������       �                      @������������������������       �                     A@-      .                    �?�<ݚ�?            �F@������������������������       �        	             .@/      >                  @m@�q�q�?             >@0      1                  `@      �?             2@������������������������       �                     @2      5                   �?���Q��?
             .@3      4                  `k@�q�q�?             @������������������������       �                     �?������������������������       �                      @6      7                  `a@�q�q�?             (@������������������������       �                     @8      ;                   @և���X�?             @9      :                  @j@���Q��?             @������������������������       �                      @������������������������       �                     @<      =                  0f@      �?              @������������������������       �                     �?������������������������       �                     �??      D                   f@�8��8��?	             (@@      C                   �?      �?             @A      B                  �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @G      H                   �?��S���?             .@������������������������       �                     @I      J                  �e@���|���?             &@������������������������       �                     @K      N                   @      �?              @L      M                  �Z@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @r  tr  bh�h"h#K �r  h%�r  Rr	  (KMOKK�r
  hR�B�       �t@     y@     �T@     @o@     �R@     `d@      A@      a@      (@     @Y@      @      W@      @     �D@       @      @      �?              �?      @              @      �?              @      C@      @      7@      �?      3@              &@      �?       @              @      �?      @      �?                      @       @      @              @       @      �?              �?       @                      .@      �?     �I@              F@      �?      @      �?                      @      @      "@      @                      "@      6@      B@      .@      (@      @       @               @      @              (@      $@      (@      @      (@      @       @      @              @       @              $@                       @              @      @      8@      @      4@       @      4@       @      @              @       @                      0@      �?              @      @              @      @      �?      @                      �?      D@      :@      <@      :@      8@      :@      6@      1@      �?      @      �?                      @      5@      *@      @       @      @      �?              �?      @                      �?      ,@      &@      @      @       @       @              �?       @      �?       @                      �?      �?      @              @      �?      �?      �?                      �?      &@      @      �?      @      �?                      @      $@       @       @      �?      �?              �?      �?              �?      �?               @      �?      @              @      �?              �?      @               @      "@       @      �?      �?              �?      �?              �?      �?                       @      @              (@              "@     �U@      @     �U@      @      @      @              �?      @      �?      �?              �?      �?                      @      @     �T@      �?      @              @      �?               @     �S@              G@       @     �@@       @      &@      �?      �?              �?      �?              �?      $@      �?      @               @      �?      �?      �?                      �?              @              6@       @             @o@     �b@     �`@     �]@      @      9@      �?      5@      �?      @      �?      @              @      �?      �?              �?      �?                       @              ,@      @      @      �?      @      �?                      @       @              `@     @W@     �U@     �C@      O@      6@      J@      (@      &@      "@      &@      @              �?      &@       @      @               @       @       @      �?      @               @      �?       @                      �?              �?              @     �D@      @      0@              9@      @      *@              (@      @      (@                      @      $@      $@      @      $@              @      @      @      @      @      @                      @      @              @              8@      1@      @      �?      @      �?              �?      @              @              1@      0@      1@      (@       @      @              @       @      @               @       @      �?       @                      �?      .@      @       @      @              @       @              *@       @      @              "@       @      "@      �?      @              @      �?              �?      @                      �?              @     �E@      K@      *@     �A@      *@      A@      &@      A@      $@      A@      @      ,@      @      @      @              @      @              @      @      @      @                      @              @      @      4@              $@      @      $@      �?               @      $@       @      @              @       @                      @      �?               @                      �?      >@      3@      @      (@      �?               @      (@              $@       @       @      �?       @      �?                       @      �?              ;@      @      7@       @      (@       @      (@                       @      &@              @      @       @      @      �?              �?      @              @      �?       @               @      �?               @             @]@     �@@     �[@      9@     �[@      7@      1@      &@              @      1@       @      &@      �?      @              @      �?      @                      �?      @      @              @      @      @      @               @      @      �?      @               @      �?       @              �?      �?      �?      �?                      �?      �?             @W@      (@      M@       @      8@       @      8@                       @      A@             �A@      $@      .@              4@      $@      "@      "@              @      "@      @      �?       @      �?                       @       @      @      @              @      @       @      @       @                      @      �?      �?              �?      �?              &@      �?      @      �?       @      �?              �?       @              �?               @                       @      @       @              @      @      @      @              @      @      @       @               @      @                       @r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h8Kh9Kh:h"h#K �r  h%�r  Rr  (KK�r  hR�C              �?r  tr  bhFhVhAC       r  �r  Rr  hZKh[h\Kh"h#K �r  h%�r  Rr  (KK�r  hA�C       r  tr  bK�r  Rr  }r   (hKhfMhgh"h#K �r!  h%�r"  Rr#  (KM�r$  hn�B�>         �                    �?6������?�           ��@       3                   `_@d}h���?�            �w@       (                   �`@�?�P�a�?s            �f@                            �?|�H���?7            �V@                          @_@�z�G��?             $@                           ]@և���X�?             @������������������������       �                     �?                           �?      �?             @	       
                    Z@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @       '                    y@����?�?1            @T@                          h@p#�����?0            �S@                           �?��S�ۿ?            �F@                          �Z@H%u��?             9@������������������������       �                     �?                           _@�8��8��?             8@������������������������       �                     &@                           `@8�Z$���?             *@������������������������       �                      @������������������������       �                     &@������������������������       �                     4@       &                   �p@������?             A@       %                    �?�ՙ/�?             5@       $                   �o@D�n�3�?             3@                           Z@������?             .@                          �l@���Q��?             @������������������������       �                     @������������������������       �                      @        #                   @Z@ףp=
�?             $@!       "                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     *@������������������������       �                      @)       2                   �K@ }�Я��?<            @V@*       1                    �?Pa�	�?            �@@+       ,                   `]@��S�ۿ?             .@������������������������       �                     $@-       .                   @b@z�G�z�?             @������������������������       �                     @/       0                   @^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             2@������������������������       �        '             L@4       �                    �?:ɨ��?}            �h@5       D                   p`@䯦s#�?b            �c@6       C                   `p@���Q��?             9@7       8                   �h@�X����?             6@������������������������       �                     @9       @                   p`@j���� �?	             1@:       ?                    `@�	j*D�?             *@;       >                   �_@ףp=
�?             $@<       =                   0k@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @A       B                     �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @E       �                   �f@��C�?S            �`@F       U                    �?FVQ&�?Q            �`@G       T                   �c@b�h�d.�?            �A@H       O                   �[@�+e�X�?             9@I       J                   �g@�q�q�?             @������������������������       �                     �?K       L                    c@z�G�z�?             @������������������������       �                      @M       N                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @P       S                   `a@�KM�]�?             3@Q       R                   c@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     (@������������������������       �                     $@V       g                     �?@��Pl3�?=            @X@W       f                   �s@�\��N��?             3@X       c                   �c@      �?
             0@Y       \                   Pm@���!pc�?             &@Z       [                    [@      �?             @������������������������       �                      @������������������������       �                      @]       ^                   ``@؇���X�?             @������������������������       �                     @_       `                   �a@      �?             @������������������������       �                      @a       b                   `b@      �?              @������������������������       �                     �?������������������������       �                     �?d       e                   �m@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @h       q                   @g@�99lMt�?1            �S@i       j                   @Y@�q�q�?
             (@������������������������       �                     @k       l                   �`@X�<ݚ�?             "@������������������������       �                     �?m       n                   �a@      �?              @������������������������       �                     @o       p                   pf@���Q��?             @������������������������       �                     @������������������������       �                      @r       �                   �b@:ɨ��?'            �P@s       �                   0c@�BbΊ�?#             M@t       �                   �`@��2(&�?             F@u       ~                    �?�θ�?             :@v       y                   pj@�KM�]�?             3@w       x                   `i@      �?             @������������������������       �                     @������������������������       �                     �?z       {                   @_@��S�ۿ?	             .@������������������������       �                     $@|       }                   8s@z�G�z�?             @������������������������       �                     �?������������������������       �                     @       �                   �n@և���X�?             @������������������������       �                     @�       �                   pa@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             2@�       �                    b@X�Cc�?
             ,@�       �                    \@�	j*D�?	             *@�       �                   pd@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �c@z�G�z�?             $@������������������������       �                     @�       �                    a@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                   �a@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                    �C@�       �                    �?J����*�?�            @v@�       �                    _@�W���?e            @d@�       �                   �Z@tk~X��?-             R@������������������������       �                     @�       �                   �c@<���D�?*            �P@�       �                   (p@�g�y��?             ?@������������������������       �                     5@�       �                    �?ףp=
�?             $@������������������������       �                     �?�       �                   xp@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                   Pl@z�G�z�?            �A@������������������������       �                     1@�       �                   e@b�2�tk�?
             2@�       �                    �?�z�G��?             $@�       �                   r@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   �^@(;L]n�?8            �V@�       �                   �^@���!pc�?             &@�       �                   �b@z�G�z�?             $@������������������������       �                     @�       �                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �        0            �S@�       �                   P`@�-p%���?x            @h@�       �                    T@PN���?>            @V@�       �                    �?     ��?             0@�       �                    �?d}h���?	             ,@�       �                   �Z@�<ݚ�?             "@������������������������       �                     @�       �                   �\@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    @z�G�z�?             @�       �                    _@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    ]@&��f���?3            @R@�       �                    f@8�A�0��?             6@�       �                   �p@��.k���?
             1@�       �                    @      �?             (@�       �                   �[@z�G�z�?             $@�       �                   `m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �_@�t����?&            �I@�       �                    @ �q�q�?             8@�       �                    �?�X�<ݺ?             2@�       �                    �?�IєX�?             1@������������������������       �                     @�       �                   �s@$�q-�?             *@������������������������       �        	             &@�       �                     �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �o@�+$�jP�?             ;@�       �                   �j@�����?             5@������������������������       �                     "@�       �                   �j@r�q��?             (@������������������������       �                     �?�       �                   l@�C��2(�?
             &@������������������������       �                     @�       �                    `@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                     �?      �?             @�       �                   �]@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   c@�xGZ���?:            @Z@�       �                   �`@д>��C�?             =@�       �                    ]@�8��8��?             8@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             5@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �`@��}�+r�?,             S@������������������������       �                      @�                            �?` .�(�?+            �R@�       �                    @�X�<ݺ?             2@�       �                   0e@�8��8��?             (@������������������������       �                     "@�       �                   @q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                         @���>4��?              L@      	                  �`@�>$�*��?            �D@                        0b@     ��?             0@������������������������       �                     @                        �\@�q�q�?             "@������������������������       �                     @                         _@      �?             @������������������������       �                     @������������������������       �                     @
                        `a@z�G�z�?             9@������������������������       �                     &@                         �?X�Cc�?             ,@                         b@X�<ݚ�?             "@                        �n@և���X�?             @                         �?���Q��?             @                        �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                        �l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        f@z�G�z�?	             .@                        �o@؇���X�?             ,@                        �b@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?r%  tr&  bh�h"h#K �r'  h%�r(  Rr)  (KMKK�r*  hR�B�       �t@     �x@     @T@     �r@      5@     �c@      4@     �Q@      @      @      @      @      �?              @      @      �?      @              @      �?               @              @              *@      Q@      &@      Q@      @      E@      @      6@      �?               @      6@              &@       @      &@       @                      &@              4@       @      :@       @      *@       @      &@      @      &@      @       @      @                       @      �?      "@      �?      �?              �?      �?                       @      @                       @              *@       @              �?      V@      �?      @@      �?      ,@              $@      �?      @              @      �?      �?      �?                      �?              2@              L@      N@     @a@      N@     �X@      .@      $@      .@      @      @              $@      @      "@      @      "@      �?      @      �?      @                      �?      @                      @      �?      @      �?                      @              @     �F@     @V@     �E@     @V@      @      =@      @      3@      @       @              �?      @      �?       @               @      �?              �?       @               @      1@       @      @              @       @                      (@              $@     �B@      N@      "@      $@      @      $@      @       @       @       @       @                       @      �?      @              @      �?      @               @      �?      �?      �?                      �?      @       @      @                       @      @              <@      I@       @      @      @              @      @              �?      @      @      @               @      @              @       @              4@      G@      .@     �E@      @      C@      @      4@       @      1@      �?      @              @      �?              �?      ,@              $@      �?      @      �?                      @      @      @      @              �?      @      �?                      @              2@      "@      @      "@      @      �?       @      �?                       @       @       @      @              @       @      @                       @              �?      @      @      @                      @       @                     �C@     �o@     �Y@      b@      1@      M@      ,@              @      M@       @      >@      �?      5@              "@      �?      �?               @      �?              �?       @              <@      @      1@              &@      @      @      @       @      @              @       @              �?               @             �U@      @       @      @       @       @      @              �?       @      �?                       @              �?     �S@             @[@     @U@     �N@      <@      @      *@      @      &@       @      @              @       @      @       @                      @      �?      @      �?      @      �?                      @              �?               @      M@      .@      *@      "@       @      "@      @      "@       @       @       @      �?       @                      �?              @      �?      �?      �?                      �?      @              @             �F@      @      7@      �?      1@      �?      0@      �?      @              (@      �?      &@              �?      �?      �?                      �?      �?              @              6@      @      3@       @      "@              $@       @              �?      $@      �?      @              @      �?              �?      @              @      @       @       @               @       @              �?      �?              �?      �?              H@     �L@      @      8@       @      6@       @      �?       @                      �?              5@      @       @      @                       @     �E@     �@@               @     �E@      ?@      1@      �?      &@      �?      "@               @      �?              �?       @              @              :@      >@      7@      2@      @      *@              @      @      @              @      @      @      @                      @      4@      @      &@              "@      @      @      @      @      @      @       @      �?       @               @      �?               @                       @      �?      �?              �?      �?              @              @      (@       @      (@       @      @              @       @                      @      �?        r+  tr,  bubhhubh)�r-  }r.  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h8Kh9Kh:h"h#K �r/  h%�r0  Rr1  (KK�r2  hR�C              �?r3  tr4  bhFhVhAC       r5  �r6  Rr7  hZKh[h\Kh"h#K �r8  h%�r9  Rr:  (KK�r;  hA�C       r<  tr=  bK�r>  Rr?  }r@  (hKhfMhgh"h#K �rA  h%�rB  RrC  (KM�rD  hn�B=         �                    �?U�ք�?�           ��@       =                   P`@r=ά�{�?�            Px@                          Ph@��M�'�?�            �k@                           �?��<b�ƥ?5             W@������������������������       �        &             Q@                           [@�8��8��?             8@������������������������       �                     &@                           �?8�Z$���?             *@	       
                   �\@"pc�
�?             &@������������������������       �                     �?                           `@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                      @       .                   p`@HX���?Q            ``@                            �?�+e�X�?!             I@                          @_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?       !                   `_@:	��ʵ�?            �F@                            `@�FVQ&�?            �@@                          �Z@�C��2(�?             6@                           �?"pc�
�?             &@������������������������       �                     �?                          @o@ףp=
�?             $@������������������������       �                     @                           Y@z�G�z�?             @������������������������       �                      @                          �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@������������������������       �                     &@"       +                    �?      �?             (@#       *                    �?r�q��?             @$       %                   �h@z�G�z�?             @������������������������       �                      @&       )                    `@�q�q�?             @'       (                   �k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?,       -                    `@r�q��?             @������������������������       �                     @������������������������       �                     �?/       0                   0q@ 7���B�?0            @T@������������������������       �                     �I@1       6                   �]@ףp=
�?             >@2       5                    �?�}�+r��?
             3@3       4                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@7       :                    �?"pc�
�?             &@8       9                   �r@؇���X�?             @������������������������       �                     �?������������������������       �                     @;       <                    �?      �?             @������������������������       �                     �?������������������������       �                     @>       �                    �?�)��V��?m            �d@?       t                   `a@�9mf��?U            �_@@       [                   `\@��6���?9             U@A       L                   �b@���|���?            �@@B       C                   �U@��S���?             .@������������������������       �                     @D       K                   �n@�q�q�?
             (@E       F                    a@X�<ݚ�?             "@������������������������       �                     @G       H                   �a@r�q��?             @������������������������       �                     @I       J                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @M       R                    �?�<ݚ�?             2@N       Q                   �[@����X�?             @O       P                   0l@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @S       Z                   �e@"pc�
�?             &@T       U                     �?ףp=
�?             $@������������������������       �                      @V       W                   pc@      �?              @������������������������       �                     @X       Y                   pd@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?\       s                    �?�q�q�?"            �I@]       b                    _@���Q �?             �H@^       a                   �c@z�G�z�?             4@_       `                   �a@���|���?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     "@c       f                     �?П[;U��?             =@d       e                   @v@$�q-�?	             *@������������������������       �                     (@������������������������       �                     �?g       l                   0j@      �?             0@h       k                   ``@�q�q�?             @i       j                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?m       n                    `@8�Z$���?	             *@������������������������       �                     @o       r                   �`@�q�q�?             @p       q                   8s@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @u       v                   �e@����X�?             E@������������������������       �                     @w       x                    c@r�q��?             B@������������������������       �                     5@y       z                   l@���Q��?
             .@������������������������       �                     @{       |                   Po@�q�q�?             "@������������������������       �                     @}       �                    e@      �?             @~                           b@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   @l@z�G�z�?             D@������������������������       �                     5@�       �                   �b@D�n�3�?             3@�       �                   �a@z�G�z�?             $@�       �                    m@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �                     �? �>�?�            �u@�       �                    �?h�WH��?A             [@�       �                    \@@4և���?:            �X@�       �                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                   �a@@��,B�?6            �V@�       �                   pa@      �?             @@������������������������       �                     <@�       �                    �?      �?             @�       �                   p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        $            �M@�       �                   �d@�z�G��?             $@�       �                   �a@      �?              @������������������������       �                     @�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?�����?�            �m@�       �                   �e@z�09JX�??            @X@�       �                   �_@ ��~���?<            �V@�       �                   �a@z�G�z�?             D@�       �                   p@      �?              @�       �                   �[@���Q��?             @������������������������       �                     �?�       �                   �T@      �?             @������������������������       �                     �?�       �                   @j@�q�q�?             @������������������������       �                     �?�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?     ��?             @@�       �                   �\@ܷ��?��?             =@�       �                   `c@z�G�z�?             @������������������������       �                     @�       �                    f@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�8��8��?             8@�       �                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �p@���7�?             6@������������������������       �                     2@�       �                    d@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    `@ףp=
�?             I@�       �                   �^@�q�q�?             (@�       �                   @n@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     C@�       �                   `p@����X�?             @������������������������       �                      @������������������������       �                     @�       �                   �_@B� ��?Z            �a@�       �                    �?��-�=��?            �C@�       �                   Xr@�㙢�c�?             7@�       �                   @]@؇���X�?             5@�       �                   �j@z�G�z�?
             .@�       �                   �`@���!pc�?             &@������������������������       �                     @�       �                   �U@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@�       
                   �?<�;�OK�?@            @Y@�       �                   @[@��]�T��?4            �T@������������������������       �                     @�       �                    @v�_���?3            �S@�       �                    T@^(��I�?&            �K@�       �                    d@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   pg@H.�!���?#             I@������������������������       �                      @�       �                   `a@0,Tg��?             E@�       �                   p`@���y4F�?             C@�       �                   �j@r٣����?            �@@�       �                   �g@�q�q�?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                   �b@PN��T'�?             ;@������������������������       �                     $@�       �                    �?������?             1@�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    ]@d}h���?             ,@�       �                    f@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �b@r�q��?             (@������������������������       �                      @������������������������       �                     $@������������������������       �                     @�       �                    �?      �?             @�       �                   `d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @       	                   p@r�q��?             8@                        b@b�2�tk�?	             2@������������������������       �                      @                        @_@�z�G��?             $@������������������������       �                      @                        0f@      �?              @������������������������       �                     @                         a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                         �?�����?             3@                        0o@������?
             1@                         �?      �?              @                        @]@�q�q�?             @������������������������       �                     �?������������������������       �                      @                        �a@���Q��?             @                        �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     "@������������������������       �                      @rE  trF  bh�h"h#K �rG  h%�rH  RrI  (KMKK�rJ  hR�Bp        t@     �y@     �T@      s@      1@     �i@       @     �V@              Q@       @      6@              &@       @      &@       @      "@      �?              �?      "@      �?                      "@               @      .@      ]@      (@      C@      @      �?      @                      �?       @     �B@       @      ?@       @      4@       @      "@      �?              �?      "@              @      �?      @               @      �?       @               @      �?                      &@              &@      @      @      �?      @      �?      @               @      �?       @      �?      �?      �?                      �?              �?              �?      @      �?      @                      �?      @     �S@             �I@      @      ;@      �?      2@      �?      @              @      �?                      &@       @      "@      �?      @      �?                      @      �?      @      �?                      @     �P@      Y@      M@      Q@      G@      C@      (@      5@       @      @      @              @      @      @      @              @      @      �?      @               @      �?       @                      �?              @      @      ,@       @      @       @      @              @       @                       @       @      "@      �?      "@               @      �?      @              @      �?      @      �?                      @      �?              A@      1@      @@      1@      0@      @      @      @      @                      @      "@              0@      *@      (@      �?      (@                      �?      @      (@       @      �?      �?      �?              �?      �?              �?               @      &@              @       @      @       @       @       @                       @               @       @              (@      >@      @              @      >@              5@      @      "@              @      @      @      @              @      @      �?      @      �?                      @       @               @      @@              5@       @      &@       @       @      @       @      @                       @      @                      "@     �m@     �Z@     �X@      $@     �V@      @      �?      @              @      �?             �V@      �?      ?@      �?      <@              @      �?      �?      �?      �?                      �?       @             �M@              @      @      @      �?      @               @      �?              �?       @                       @     �a@      X@     �S@      2@     @S@      *@      @@       @      @      @      @       @      �?               @       @              �?       @      �?      �?              �?      �?              �?      �?                      @      =@      @      :@      @      @      �?      @              �?      �?              �?      �?              6@       @      �?      �?              �?      �?              5@      �?      2@              @      �?              �?      @              @             �F@      @      @      @      @      �?      @                      �?              @      C@               @      @       @                      @      O@     �S@      @     �A@      @      3@      @      2@      @      (@      @       @              @      @      �?              �?      @                      @              @      �?      �?              �?      �?                      0@      M@     �E@      J@      >@              @      J@      ;@     �D@      ,@       @      @       @                      @     �C@      &@       @              ?@      &@      >@       @      9@       @       @      @               @       @       @       @                       @      7@      @      $@              *@      @       @      �?              �?       @              &@      @      �?      �?              �?      �?              $@       @               @      $@              @              �?      @      �?      �?              �?      �?                       @      &@      *@      &@      @       @              @      @       @              �?      @              @      �?       @               @      �?                      @      @      *@      @      *@      @      @       @      �?              �?       @               @      @       @      �?              �?       @                       @              "@       @        rK  trL  bubhhubh)�rM  }rN  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h8Kh9Kh:h"h#K �rO  h%�rP  RrQ  (KK�rR  hR�C              �?rS  trT  bhFhVhAC       rU  �rV  RrW  hZKh[h\Kh"h#K �rX  h%�rY  RrZ  (KK�r[  hA�C       r\  tr]  bK�r^  Rr_  }r`  (hKhfMChgh"h#K �ra  h%�rb  Rrc  (KMC�rd  hn�B�F         6                     �?0����?�           ��@       /                    �?�-١�:�?]            @a@                           a@�p�I�?Q            �]@                           �?Du9iH��?8            �U@                           �?"pc�
�?             6@������������������������       �                     @                          �i@������?             1@       	                   @[@      �?             @������������������������       �                      @
                           `@      �?             @������������������������       �                     @������������������������       �                     �?                           �?�C��2(�?             &@                          �p@؇���X�?             @������������������������       �                     @                          �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          �Z@      �?*             P@                           �?�q�q�?             @                           @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �        '            �N@       .                   8s@�'�=z��?            �@@       %                   �b@և���X�?             <@                           �]@@�0�!��?             1@                          @o@      �?             @������������������������       �                      @������������������������       �                      @!       "                   �a@$�q-�?	             *@������������������������       �                     @#       $                   �a@؇���X�?             @������������������������       �                     �?������������������������       �                     @&       -                   �r@"pc�
�?	             &@'       ,                    d@ףp=
�?             $@(       )                   `a@z�G�z�?             @������������������������       �                      @*       +                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @0       5                    �?�����?             3@1       4                   �p@և���X�?	             ,@2       3                   �]@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @7       �                    �?��Vu@z�?y           ��@8       �                   @d@X���o�?�            �u@9       �                    �?*)��?�            �t@:       _                   `_@����o�?�            �o@;       >                   �Z@4Qi0���?I            �^@<       =                    ]@�q�q�?             @������������������������       �                      @������������������������       �                     �??       R                   �`@��(\���?F             ^@@       C                    V@�����H�?              K@A       B                    �?���Q��?             @������������������������       �                     @������������������������       �                      @D       K                    �?Hm_!'1�?            �H@E       J                    I@��Y��]�?            �D@F       G                   �Z@�����H�?             "@������������������������       �                     @H       I                   �[@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @@L       M                   �^@      �?              @������������������������       �                     @N       Q                   �Y@���Q��?             @O       P                    `@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @S       T                   �Z@���7�?&            �P@������������������������       �                     9@U       ^                   �l@��p\�?            �D@V       Y                   �[@      �?             8@W       X                   �b@      �?             @������������������������       �                      @������������������������       �                      @Z       [                   �b@P���Q�?             4@������������������������       �                     2@\       ]                   @^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             1@`       �                   �b@�G\�c�?O            @`@a       �                   �e@d}h��?F             \@b       �                   `o@���vq�?C            �Z@c       z                   �k@���Q��?,            @P@d       e                   `@�q�q�?             E@������������������������       �                     @f       y                    �?�d�����?             C@g       j                    �?     ��?             @@h       i                   �i@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @k       v                   �`@�LQ�1	�?             7@l       u                   pj@j���� �?             1@m       n                   �a@��
ц��?
             *@������������������������       �                     @o       t                   @_@���Q��?             $@p       s                   �\@      �?              @q       r                   pc@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @w       x                   �g@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @{       �                   �a@
;&����?             7@|       }                   l@և���X�?             5@������������������������       �                     @~                          �`@��.k���?             1@������������������������       �                     @�       �                   �m@�q�q�?	             (@�       �                   �m@և���X�?             @�       �                   �b@      �?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �a@��r._�?            �D@�       �                   `a@�z�G��?
             4@������������������������       �                     $@�       �                   �p@���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                   0c@���N8�?             5@������������������������       �                     $@�       �                   `q@�C��2(�?             &@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   P`@r�q��?	             2@������������������������       �                      @�       �                    �?      �?             0@�       �                    f@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   s@ �\���?0            �S@�       �                   @a@ �й���?,            @R@������������������������       �                    �H@�       �                   �^@ �q�q�?             8@������������������������       �        	             (@�       �                    �?�8��8��?             (@�       �                   @a@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   `t@      �?             @������������������������       �                     �?�       �                    y@���Q��?             @������������������������       �                      @�       �                   ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �p@�}�+r��?             3@������������������������       �        	             *@�       �                    �?r�q��?             @������������������������       �                      @�       �                   �q@      �?             @������������������������       �                     �?������������������������       �                     @�       .                   �?f���?�            �n@�       #                   @����X�?�            `i@�       �                   @\@���"͏�?z             g@�       �                   @Y@b�2�tk�?             2@�       �                   `X@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?      �?             (@�       �                    �?�q�q�?             "@������������������������       �                      @�       �                   @[@և���X�?             @������������������������       �                      @�       �                   @^@���Q��?             @������������������������       �                      @�       �                   `_@�q�q�?             @������������������������       �                     �?�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    ]@$Z9��?m            �d@�       �                    �?�G��l��?             5@�       �                   pf@      �?             4@�       �                    Z@      �?             0@������������������������       �                      @�       �                   �k@և���X�?             ,@������������������������       �                     @�       �                    �?z�G�z�?             $@������������������������       �                     @�       �                   �Z@�q�q�?             @������������������������       �                     �?�       �                   @[@z�G�z�?             @������������������������       �                      @�       �                   �p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?�@i����?]            @b@�       �                   0d@r֛w���?             ?@�       �                    b@p�ݯ��?             3@�       �                    Z@      �?              @�       �                   Pb@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �b@�eP*L��?             &@������������������������       �                     @�       �                   0c@����X�?             @������������������������       �                     @�       �                    `@�q�q�?             @������������������������       �                     �?�       �                   �k@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    e@�8��8��?	             (@������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     @�       �                   q@      �?              @������������������������       �                     �?������������������������       �                     �?�                          �?�LQ�1	�?H            �\@�       �                   Hp@�.ߴ#�?(            �N@������������������������       �                    �B@�                          d@      �?             8@�                          �_@�θ�?             *@������������������������       �                      @                        �a@�C��2(�?             &@������������������������       �                     @                        �q@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@      "                  c@�<ݚ�?              K@                        0d@���B���?             J@	                         T@      �?              @
                        �^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                        �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        `a@�C��2(�?             F@                        �g@��S�ۿ?             >@                        �f@      �?              @������������������������       �                     �?������������������������       �                     �?                        �b@h�����?             <@                        @_@��S�ۿ?	             .@                        0m@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@      !                  �d@؇���X�?             ,@                        �a@      �?              @������������������������       �                     @                          �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @$      -                   �?�E��ӭ�?             2@%      (                  0`@�n_Y�K�?	             *@&      '                  �m@      �?             @������������������������       �                     @������������������������       �                     �?)      *                  �d@�<ݚ�?             "@������������������������       �                     @+      ,                  �c@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @/      @                  �j@և���X�?             E@0      5                  �_@�'�=z��?            �@@1      4                   �?�r����?             .@2      3                  �i@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     "@6      ;                   j@r�q��?             2@7      8                   �?@4և���?
             ,@������������������������       �                     @9      :                  @e@�����H�?             "@������������������������       �                      @������������������������       �                     �?<      ?                   �?      �?             @=      >                  �j@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?A      B                  �c@�����H�?             "@������������������������       �                      @������������������������       �                     �?re  trf  bh�h"h#K �rg  h%�rh  Rri  (KMCKK�rj  hR�B0        u@     �x@     �Y@     �A@     @X@      6@      T@      @      2@      @      @              *@      @      @      @       @              �?      @              @      �?              $@      �?      @      �?      @              �?      �?      �?                      �?      @              O@       @      �?       @      �?      �?              �?      �?                      �?     �N@              1@      0@      (@      0@      @      ,@       @       @       @                       @      �?      (@              @      �?      @      �?                      @      "@       @      "@      �?      @      �?       @               @      �?       @                      �?      @                      �?      @              @      *@      @       @       @       @       @                       @      @                      @      m@     �v@     �Q@     �q@     @Q@     pp@     @P@     �g@      &@      \@       @      �?       @                      �?      "@     �[@      @      H@       @      @              @       @              @     �F@      �?      D@      �?       @              @      �?      @      �?                      @              @@      @      @              @      @       @      �?       @      �?                       @       @              @     �O@              9@      @      C@      @      5@       @       @       @                       @      �?      3@              2@      �?      �?      �?                      �?              1@      K@      S@     �C@     @R@     �@@     @R@      :@     �C@      ,@      <@      @              $@      <@      $@      6@       @      @              @       @               @      .@      @      $@      @      @      @              @      @       @      @       @      @              @       @                      @       @                      @      �?      @      �?                      @              @      (@      &@      (@      "@      @               @      "@              @       @      @      @      @      @      �?       @      �?              �?       @              �?              �?       @               @      �?              @      �?              �?      @                       @      @      A@      @      ,@              $@      @      @              @      @              �?      4@              $@      �?      $@      �?       @              �?      �?      �?              �?      �?                       @      @              .@      @               @      .@      �?       @      �?       @                      �?      @              @     �R@      �?      R@             �H@      �?      7@              (@      �?      &@      �?      @              @      �?                      @      @      @      �?               @      @               @       @      �?       @                      �?      �?      2@              *@      �?      @               @      �?      @      �?                      @     `d@     �T@      b@      M@     �a@     �F@      @      &@      @       @               @      @              @      "@      @      @               @      @      @               @      @       @       @              �?       @              �?      �?      �?      �?                      �?              @     �`@      A@      $@      &@      $@      $@      @      $@               @      @       @      @               @       @              @       @      @      �?              �?      @               @      �?       @               @      �?              @                      �?     �^@      7@      7@       @      (@      @      @      �?      �?      �?              �?      �?              @              @      @              @      @       @      @              �?       @              �?      �?      �?              �?      �?              &@      �?      @              @      �?      @              �?      �?              �?      �?              Y@      .@      M@      @     �B@              5@      @      $@      @               @      $@      �?      @              @      �?      @                      �?      &@              E@      (@      E@      $@       @      @      �?      @      �?                      @      �?       @               @      �?              D@      @      <@       @      �?      �?      �?                      �?      ;@      �?      ,@      �?      @      �?      @                      �?       @              *@              (@       @      @       @      @              �?       @               @      �?              @                       @      @      *@      @       @      @      �?      @                      �?       @      @              @       @      @       @                      @              @      2@      8@      1@      0@       @      *@       @      @              @       @                      "@      .@      @      *@      �?      @               @      �?       @                      �?       @       @      �?       @               @      �?              �?              �?       @               @      �?        rk  trl  bubhhubh)�rm  }rn  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h8Kh9Kh:h"h#K �ro  h%�rp  Rrq  (KK�rr  hR�C              �?rs  trt  bhFhVhAC       ru  �rv  Rrw  hZKh[h\Kh"h#K �rx  h%�ry  Rrz  (KK�r{  hA�C       r|  tr}  bK�r~  Rr  }r�  (hKhfM+hgh"h#K �r�  h%�r�  Rr�  (KM+�r�  hn�BhA         �                   �`@�+	G�?�           ��@       k                    �?l�"�^%�?�            �u@       <                    �?0�	B��?�            �n@                          �h@h�_���?q            `e@                           _@
��[��?(            @P@                          �g@r�����?            �J@                          �b@>a�����?            �I@       	                   �Z@�*/�8V�?            �G@������������������������       �        	             ,@
                           I@6YE�t�?            �@@                           `@�d�����?             3@                          `\@����X�?             @������������������������       �                     @                           �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     (@������������������������       �                     ,@                          @c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                          �Y@�q�q�?	             (@������������������������       �                      @                          @d@z�G�z�?             $@                          `_@�����H�?             "@                          0a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?        )                     �?�8�l��?I            �Z@!       (                   �`@8�Z$���?	             *@"       %                    �?�q�q�?             @#       $                   �k@      �?             @������������������������       �                     @������������������������       �                     �?&       '                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @*       3                   �k@ rpa�?@            @W@+       ,                    �?�r����?             >@������������������������       �                     4@-       .                   �\@���Q��?             $@������������������������       �                      @/       0                   @_@      �?              @������������������������       �                     @1       2                   �k@���Q��?             @������������������������       �                     @������������������������       �                      @4       ;                   `\@ ������?,            �O@5       :                   pp@�nkK�?             7@6       9                   �`@؇���X�?             @7       8                   o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     0@������������������������       �                     D@=       R                    \@p�ݯ��?1             S@>       C                   �V@�q�q�?             8@?       @                    �?      �?             @������������������������       �                      @A       B                   @\@      �?              @������������������������       �                     �?������������������������       �                     �?D       Q                    �?      �?             4@E       H                     �?�n_Y�K�?	             *@F       G                    @���Q��?             @������������������������       �                     @������������������������       �                      @I       J                    W@      �?              @������������������������       �                     @K       L                   �X@���Q��?             @������������������������       �                     �?M       N                    �?      �?             @������������������������       �                      @O       P                    Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @S       T                    �?�θ�?"             J@������������������������       �        	             .@U       Z                   @]@4�B��?            �B@V       Y                   �\@�����H�?             "@W       X                    ]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @[       \                   �]@��>4և�?             <@������������������������       �                      @]       ^                   �c@$��m��?             :@������������������������       �                     @_       j                   �a@�GN�z�?             6@`       i                    �?�q�q�?	             .@a       b                     �?����X�?             ,@������������������������       �                      @c       f                    @�q�q�?             (@d       e                   �`@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @g       h                   `]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @l       m                   ``@�C��2(�?A            �X@������������������������       �                     A@n       o                   �k@��ɉ�?)            @P@������������������������       �                     @@p       q                   �`@���!pc�?            �@@������������������������       �                     �?r       s                   �[@      �?             @@������������������������       �                      @t                           �?�q�q�?             8@u       v                   Pa@�n_Y�K�?             *@������������������������       �                     @w       z                   �]@z�G�z�?             $@x       y                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?{       |                   �a@      �?              @������������������������       �                     @}       ~                   �o@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@�                         �a@�E���?�            @x@�       �                    �?�/� ��?�            �s@�       �                    �?�����?�             q@�       �                     �?�ҿf���?2            �T@�       �                    �?D�n�3�?             3@������������������������       �                     @�       �                    �?      �?             0@�       �                   �\@�n_Y�K�?             *@������������������������       �                     @�       �                   �q@����X�?             @������������������������       �                     @�       �                   c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �^@     8�?'             P@�       �                    �?�g�y��?             ?@�       �                    �?��
ц��?             :@�       �                    ]@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   pc@      �?             6@�       �                   �_@X�Cc�?	             ,@������������������������       �                      @�       �                   �a@      �?             (@�       �                   �p@      �?              @�       �                   �\@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    \@      �?              @�       �                   pi@���Q��?             @������������������������       �                     �?�       �                   �d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �n@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �l@�q�q�?            �@@�       �                   �_@      �?	             0@������������������������       �                      @�       �                   0a@؇���X�?             ,@������������������������       �                     @�       �                   0c@"pc�
�?             &@�       �                   `h@      �?              @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   ``@��.k���?
             1@������������������������       �                     @�       �                   �q@"pc�
�?             &@�       �                   �m@ףp=
�?             $@�       �                   0a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                     �?B�#-g�?u            �g@������������������������       �        #             N@�       �                   �c@�,A7H�?R            ``@������������������������       �                     @�       �                   �d@     ��?O             `@�       �                   pd@���j��?7             W@�       �                   pa@�������?5            �U@�       �                    @��W��?-            @R@�       �                   �a@�� =[�?*             Q@�       �                   Pa@�t����?             1@������������������������       �                     "@�       �                   �i@      �?              @�       �                   pa@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�t����?            �I@�       �                   �c@؇���X�?             <@������������������������       �                     1@�       �                   �o@���|���?             &@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?���}<S�?             7@������������������������       �                     @�       �                   �`@�t����?             1@�       �                   0n@      �?             0@������������������������       �                     *@�       �                   �b@�q�q�?             @������������������������       �                     �?�       �                   @[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   �_@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?��
ц��?             *@�       �                   pb@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �`@      �?              @������������������������       �                      @������������������������       �                     @�       �                   `m@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�X�<ݺ?             B@������������������������       �                     1@�       �                    f@�KM�]�?             3@�       �                   �e@�<ݚ�?             "@�       �                   �e@      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     $@�       �                   `]@X�<ݚ�?            �F@������������������������       �                      @�       �                   `_@��%��?            �B@������������������������       �                     @�                         Pa@`՟�G��?             ?@�                          �?��>4և�?             <@                         ``@��S�ۿ?             .@������������������������       �                     $@                        �`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @      
                    �?�θ�?             *@                        �d@z�G�z�?             @������������������������       �                     @      	                  @q@      �?              @������������������������       �                     �?������������������������       �                     �?                         @      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @                         �p@bKv���?+            @Q@                         �?��+��?            �B@                         T@��s����?             5@������������������������       �                     @                          �?������?
             .@������������������������       �                      @                         f@և���X�?             @                        �b@�q�q�?             @������������������������       �                     �?                        �f@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                        �c@      �?             0@                        �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             *@!      *                   @      �?             @@"      )                    �?��a�n`�?             ?@#      $                  �b@      �?             ,@������������������������       �                     @%      (                   �?�z�G��?             $@&      '                  8r@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     1@������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM+KK�r�  hR�B�       `t@     �y@     �T@     �p@     @R@     �e@      9@     @b@      2@     �G@      $@     �E@       @     �E@      @      E@              ,@      @      <@      @      ,@      @       @      @               @       @               @       @                      (@              ,@      @      �?      @                      �?       @               @      @               @       @       @       @      �?      �?      �?              �?      �?              @                      �?      @     �X@       @      &@       @      @      �?      @              @      �?              �?      �?      �?                      �?              @      @      V@      @      :@              4@      @      @       @               @      @              @       @      @              @       @              �?      O@      �?      6@      �?      @      �?      �?              �?      �?                      @              0@              D@      H@      <@       @      0@      @      �?       @              �?      �?      �?                      �?      @      .@      @       @       @      @              @       @              @      @              @      @       @              �?      @      �?       @              �?      �?      �?                      �?              @      D@      (@      .@              9@      (@       @      �?      @      �?              �?      @              @              1@      &@               @      1@      "@              @      1@      @      $@      @      $@      @       @               @      @      @       @      @                       @      �?       @               @      �?                      �?      @              "@     �V@              A@      "@      L@              @@      "@      8@      �?               @      8@               @       @      0@       @      @              @       @       @      �?      �?      �?                      �?      @      �?      @               @      �?       @                      �?              &@     �n@      b@     @k@     @Y@     �h@      S@      C@     �F@      &@       @      @               @       @      @       @              @      @       @      @              �?       @               @      �?              @              ;@     �B@      0@      .@      (@      ,@      �?      @              @      �?              &@      &@      @      "@       @              @      "@      @      @      �?      @      �?                      @       @                      @      @       @      @       @              �?      @      �?      @                      �?      @              @      �?      @                      �?      &@      6@       @      ,@               @       @      (@              @       @      "@       @      @       @      �?       @                      �?              @              @      "@       @              @      "@       @      "@      �?      �?      �?      �?                      �?       @                      �?      d@      ?@      N@              Y@      ?@              @      Y@      <@     �P@      :@     @P@      5@     �M@      ,@     �L@      &@      (@      @      "@              @      @      @      �?              �?      @                      @     �F@      @      8@      @      1@              @      @      @               @      @              @       @              5@       @      @              .@       @      .@      �?      *@               @      �?      �?              �?      �?              �?      �?                      �?       @      @       @                      @      @      @      @      �?              �?      @               @      @       @                      @      �?      @              @      �?              A@       @      1@              1@       @      @       @      @      �?      @               @      �?              �?       @                      �?      $@              4@      9@               @      4@      1@      @              ,@      1@      &@      1@      �?      ,@              $@      �?      @      �?                      @      $@      @      @      �?      @              �?      �?              �?      �?              @       @      @                       @      @              :@     �E@      2@      3@      @      1@              @      @      &@               @      @      @      @       @              �?      @      �?      @                      �?              �?      ,@       @      �?       @               @      �?              *@               @      8@      @      8@      @      @              @      @      @      �?      @      �?                      @      @                      1@      �?        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfM_hgh"h#K �r�  h%�r�  Rr�  (KM_�r�  hn�B�L         4                  0c@6������?�           ��@       �                    �?|��?���?�           @�@                          �U@ޭ�W[��?�            @t@������������������������       �                      @       `                   ``@2�J��?�             t@       /                    j@��ջ�A�?�             j@       .                    �?      �?B             Z@       -                   �f@^l��[B�?%             M@	       "                   �c@����>4�?$             L@
       !                   0a@�z�G��?             >@                           @Y@�c�Α�?             =@                          @E@�	j*D�?             :@                          �Z@      �?             8@������������������������       �                     �?                            �?��<b���?             7@������������������������       �                     �?                          `_@�GN�z�?             6@                          `]@�8��8��?             (@������������������������       �                     @                          �_@؇���X�?             @������������������������       �                     @������������������������       �                     �?                           �?���Q��?             $@������������������������       �                      @                           �?      �?              @                          �Z@      �?             @������������������������       �                      @������������������������       �                      @                           `@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?#       (                    �?$�q-�?             :@$       %                   `g@z�G�z�?             @������������������������       �                     @&       '                   Pa@      �?              @������������������������       �                     �?������������������������       �                     �?)       *                    `@���N8�?             5@������������������������       �                     3@+       ,                     �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     G@0       U                   �p@R�}e�.�?D             Z@1       J                   �a@�n_Y�K�?+            @P@2       ;                   �m@���j��?             G@3       :                    �?�8��8��?             8@4       9                   `@ףp=
�?             4@5       8                   �_@      �?              @6       7                   �k@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     (@������������������������       �                     @<       =                     �?      �?             6@������������������������       �                     @>       ?                   �X@     ��?             0@������������������������       �                     �?@       C                   0n@�q�q�?
             .@A       B                   �`@      �?             @������������������������       �                     �?������������������������       �                     @D       I                    �?"pc�
�?             &@E       F                   �^@�<ݚ�?             "@������������������������       �                     @G       H                   @]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @K       R                   �^@p�ݯ��?             3@L       M                   n@8�Z$���?             *@������������������������       �                     "@N       Q                    \@      �?             @O       P                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?S       T                   8p@r�q��?             @������������������������       �                     @������������������������       �                     �?V       [                    ^@$�q-�?            �C@W       X                   8r@8�Z$���?             *@������������������������       �                     "@Y       Z                     �?      �?             @������������������������       �                      @������������������������       �                      @\       ]                   �u@ ��WV�?             :@������������������������       �                     6@^       _                   �{@      �?             @������������������������       �                     �?������������������������       �                     @a       j                   �`@p9W��S�?N            �\@b       i                    �?      �?              @c       h                    �?؇���X�?             @d       e                     �?r�q��?             @������������������������       �                      @f       g                   �q@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?k       �                    �?�c�����?I            �Z@l       �                   �b@�P�����?8             U@m       t                     �?������?&            �I@n       o                   �b@���Q��?             @������������������������       �                      @p       q                   �o@�q�q�?             @������������������������       �                     �?r       s                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?u       �                   Xq@��<b���?!             G@v       �                   `b@����X�?            �A@w       x                   �d@8�Z$���?             :@������������������������       �                     "@y       �                   �a@������?             1@z       �                    �?���|���?             &@{       |                   �[@X�<ݚ�?             "@������������������������       �                     �?}       ~                    ^@      �?              @������������������������       �                      @       �                   Pi@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   �k@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     &@�       �                    �?����e��?            �@@�       �                    `@l��
I��?             ;@������������������������       �                     "@�       �                   �a@X�<ݚ�?             2@�       �                     �?����X�?             @�       �                   Xs@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   pd@���!pc�?             &@������������������������       �                     @�       �                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �Z@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    _@���7�?             6@������������������������       �                     ,@�       �                   `_@      �?              @�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �`@���R�?�            @t@�       �                    \@��ӭ�a�?2             R@�       �                    @"pc�
�?             6@�       �                   �V@؇���X�?             5@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�KM�]�?             3@�       �                    �?؇���X�?
             ,@�       �                    �?z�G�z�?             $@�       �                    �?      �?             @������������������������       �                     �?�       �                    W@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                     �?z�):���?"             I@������������������������       �                     &@�       �                    �?�e����?            �C@�       �                    @��
ц��?             :@�       �                    �?�û��|�?             7@�       �                   �\@�E��ӭ�?             2@������������������������       �                     �?�       �                    �?������?             1@�       �                   0a@      �?             @������������������������       �                      @������������������������       �                      @�       �                   `T@8�Z$���?	             *@�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �a@�C��2(�?             &@�       �                    �?r�q��?             @������������������������       �                     �?�       �                   �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?8�Z$���?	             *@�       �                   @^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@�       %                   @��cy�k�?�            �o@�                          �?X�;�^o�?�            �k@�       	                  pd@��H���?�             h@�       �                   �c@��t��?N            �\@�       �                    �?�ʈD��?<            �U@�       �                   p@t��ճC�?             F@������������������������       �                     >@�       �                   Pa@d}h���?             ,@������������������������       �                     @�       �                   0b@�q�q�?             "@������������������������       �                     �?�       �                   �r@      �?              @������������������������       �                      @������������������������       �                     @�       �                   �b@���H��?             E@�       �                   pa@������?            �D@������������������������       �        
             0@�       �                    �?�J�4�?             9@�       �                   `a@�C��2(�?             6@�       �                     �?�X�<ݺ?             2@������������������������       �                     @�       �                   �_@$�q-�?
             *@������������������������       �                     @�       �                    `@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   0c@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   Pb@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �c@�c�Α�?             =@������������������������       �                     @�       �                    �?���B���?             :@�       �                     �?�q�q�?             "@������������������������       �                     @�       �                   0d@���Q��?             @������������������������       �                     @������������������������       �                      @�                          �?�t����?             1@�       �                   �\@�r����?             .@������������������������       �                     @�                          d@z�G�z�?	             $@�                          �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?                          �?؇���X�?             @������������������������       �                      @                         q@z�G�z�?             @                        �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @
                        �p@ ��WV�?2            �S@                        �\@     ��?)             P@                        �[@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        $             M@                        �e@؇���X�?	             ,@������������������������       �                     $@                        `]@      �?             @������������������������       �                      @������������������������       �                      @                        0b@�q�q�?             ;@                        `]@�q�q�?             (@������������������������       �                     @                         �?����X�?             @������������������������       �                     @������������������������       �                      @                         V@�r����?
             .@������������������������       �                     �?                         �?@4և���?	             ,@������������������������       �                     @                         �d@      �?              @������������������������       �                     @!      "                   �?�q�q�?             @������������������������       �                     �?#      $                  @q@      �?              @������������������������       �                     �?������������������������       �                     �?&      3                   �?     ��?             @@'      .                  `l@���>4��?             <@(      )                  �a@ҳ�wY;�?	             1@������������������������       �                     @*      +                  �c@�eP*L��?             &@������������������������       �                     @,      -                  0i@����X�?             @������������������������       �                     @������������������������       �                      @/      0                  �`@"pc�
�?             &@������������������������       �                     �?1      2                   b@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @5      X                   @ι�~��?7            �U@6      Q                  �b@�7�QJW�?3            �R@7      N                   g@��a�n`�?+             O@8      E                   �?��ϭ�*�?'             M@9      :                   q@�}�+r��?             C@������������������������       �                     8@;      B                  @e@؇���X�?	             ,@<      =                   �?�C��2(�?             &@������������������������       �                     @>      A                   �?      �?             @?      @                  �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @C      D                  �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @F      M                   �?R���Q�?             4@G      L                   �?���!pc�?             &@H      K                  @_@      �?             @I      J                  pl@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     "@O      P                   �?      �?             @������������������������       �                     @������������������������       �                     �?R      U                   �?��
ц��?             *@S      T                   �?r�q��?             @������������������������       �                     @������������������������       �                     �?V      W                   e@؇���X�?             @������������������������       �                     @������������������������       �                     �?Y      Z                    �?�C��2(�?             &@������������������������       �                     @[      \                  �d@؇���X�?             @������������������������       �                      @]      ^                  p@z�G�z�?             @������������������������       �                     @������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM_KK�r�  hR�B�       �t@     �x@     �s@      u@      S@      o@       @             �R@      o@     �D@     �d@      *@     �V@      *@     �F@      &@     �F@      "@      5@       @      5@       @      2@      @      2@      �?              @      2@              �?      @      1@      �?      &@              @      �?      @              @      �?              @      @               @      @      @       @       @               @       @               @       @       @                       @       @                      @      �?               @      8@      �?      @              @      �?      �?      �?                      �?      �?      4@              3@      �?      �?      �?                      �?       @                      G@      <@      S@      9@      D@      *@     �@@       @      6@       @      2@       @      @      �?      @      �?                      @      �?                      (@              @      &@      &@      @              @      &@              �?      @      $@      @      �?              �?      @               @      "@       @      @              @       @      �?       @                      �?               @      (@      @      &@       @      "@               @       @      �?       @               @      �?              �?              �?      @              @      �?              @      B@       @      &@              "@       @       @       @                       @      �?      9@              6@      �?      @      �?                      @     �@@     @T@      @      �?      @      �?      @      �?       @              @      �?      @                      �?      �?              �?              :@      T@      9@     �M@      (@     �C@       @      @               @       @      �?      �?              �?      �?      �?                      �?      $@      B@      $@      9@      @      6@              "@      @      *@      @      @      @      @      �?              @      @               @      @      @      @                      @               @              @      @      @              @      @                      &@      *@      4@       @      3@              "@       @      $@      @       @      @      �?      @                      �?              �?      @       @              @      @       @      @                       @      @      �?              �?      @              �?      5@              ,@      �?      @      �?      �?      �?                      �?              @     �m@      V@      ?@     �D@      @      2@      @      2@      �?      �?      �?                      �?       @      1@       @      (@       @       @       @       @              �?       @      �?              �?       @                      @              @              @      �?              ;@      7@      &@              0@      7@      ,@      (@      ,@      "@      *@      @              �?      *@      @       @       @               @       @              &@       @      �?      �?              �?      �?              $@      �?      @      �?      �?              @      �?      @                      �?      @              �?      @      �?                      @              @       @      &@       @       @               @       @                      "@     �i@     �G@      h@      <@     �e@      3@     �X@      0@     �S@       @     �D@      @      >@              &@      @      @              @      @              �?      @       @               @      @             �B@      @     �B@      @      0@              5@      @      4@       @      1@      �?      @              (@      �?      @              @      �?              �?      @              @      �?      @                      �?      �?       @               @      �?                      �?      5@       @              @      5@      @      @      @      @               @      @              @       @              .@       @      *@       @      @               @       @       @      �?       @                      �?      @      �?       @              @      �?      �?      �?      �?                      �?      @               @             �R@      @     �O@      �?      @      �?      @                      �?      M@              (@       @      $@               @       @               @       @              2@      "@      @      @              @      @       @      @                       @      *@       @              �?      *@      �?      @              @      �?      @               @      �?      �?              �?      �?              �?      �?              *@      3@      *@      .@      &@      @      @              @      @              @      @       @      @                       @       @      "@      �?              �?      "@              "@      �?                      @      7@     �O@      *@      O@      @      L@      @     �J@       @      B@              8@       @      (@      �?      $@              @      �?      @      �?      �?              �?      �?                       @      �?       @      �?                       @      @      1@      @       @      @      @      �?      @      �?                      @       @                      @              "@      �?      @              @      �?              @      @      �?      @              @      �?              @      �?      @                      �?      $@      �?      @              @      �?       @              @      �?      @                      �?r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJQY%hG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfMahgh"h#K �r�  h%�r�  Rr�  (KMa�r�  hn�B8M         2                   �`@�Z���?�           ��@       1                   �e@8F�V�?c            `b@       &                    �?��1���?b             b@                           �?&�a2o��?.            @Q@                           �?fP*L��?             F@������������������������       �                     @                           �?z�G�z�?             D@                           W@�㙢�c�?             7@	       
                     �?�<ݚ�?             2@������������������������       �                      @                          @E@      �?             0@                          �`@z�G�z�?             .@                          �_@$�q-�?             *@������������������������       �                     @                          p`@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                          `b@@�0�!��?
             1@                           \@��S�ۿ?	             .@������������������������       �                     �?������������������������       �                     ,@������������������������       �                      @       %                   pb@��H�}�?             9@                          �Z@      �?             2@������������������������       �                     @                          `\@���Q��?
             .@������������������������       �                     @       $                   �a@      �?             (@        !                   P`@ףp=
�?             $@������������������������       �                     @"       #                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @'       (                     �?P�Lt�<�?4             S@������������������������       �                     @)       *                    �?��.N"Ҭ?0            @Q@������������������������       �                     E@+       0                   p`@�>����?             ;@,       -                    `@r�q��?
             (@������������������������       �                      @.       /                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     .@������������������������       �                      @3       �                   �`@�)����?x           X�@4       Q                     �?�2��?�            �m@5       N                    �?�5��
J�?             G@6       ?                   @l@�eP*L��?             6@7       8                    �?�q�q�?             "@������������������������       �                      @9       :                   �[@և���X�?             @������������������������       �                     @;       <                    f@      �?             @������������������������       �                      @=       >                    _@      �?              @������������������������       �                     �?������������������������       �                     �?@       K                    �?�	j*D�?             *@A       F                    ]@���!pc�?             &@B       E                   �Z@؇���X�?             @C       D                    p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @G       H                   �_@      �?             @������������������������       �                     �?I       J                   Xs@�q�q�?             @������������������������       �                      @������������������������       �                     �?L       M                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?O       P                   @e@ �q�q�?             8@������������������������       �                     7@������������������������       �                     �?R       U                   �U@�_�.��?|            �g@S       T                   @b@      �?              @������������������������       �                     @������������������������       �                      @V       ]                   �X@
aJ���?v            �f@W       X                   �W@`2U0*��?             9@������������������������       �                     (@Y       Z                    �?$�q-�?             *@������������������������       �                     $@[       \                   @^@�q�q�?             @������������������������       �                      @������������������������       �                     �?^       �                    �?̘SJl��?g            �c@_       �                   ps@t��%�?K            �\@`       a                    �?���z�k�?C            �Y@������������������������       �                     7@b       �                   8s@\���(\�?3             T@c       z                    _@�+ت�M�?2            �S@d       y                    \@��ϭ�*�?"             M@e       p                   `[@4?,R��?             B@f       o                    �?@4և���?	             ,@g       h                   �Y@ףp=
�?             $@������������������������       �                     @i       n                   �Z@؇���X�?             @j       m                   @q@r�q��?             @k       l                   �m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @q       v                    �?"pc�
�?             6@r       s                   0l@�IєX�?	             1@������������������������       �                     ,@t       u                   �n@�q�q�?             @������������������������       �                     �?������������������������       �                      @w       x                   �`@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     6@{       �                    �?���N8�?             5@|       �                   �_@�	j*D�?
             *@}       �                   `_@և���X�?             @~                           �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   a@���Q��?             @�       �                   �k@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    b@r�q��?             @�       �                   0a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �_@      �?              @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     (@�       �                    �?�+��<��?            �E@�       �                   @e@X�Cc�?             <@�       �                   `c@���Q��?             9@�       �                    �?�X����?             6@�       �                    �?؇���X�?             @�       �                   8p@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �a@���Q��?	             .@�       �                   `^@�q�q�?             "@������������������������       �                     �?�       �                   �q@      �?              @�       �                   @_@      �?             @������������������������       �                     �?�       �                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?��S�ۿ?
             .@�       �                   �]@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       :                  �a@B0�8���?�            �u@�       �                   �n@ .~�`��?�             r@�       �                    �?�IA��?g            �c@�       �                    �?|�-蝉�?Z            �`@�       �                    �?p�ݯ��?             C@�       �                     �?^������?            �A@������������������������       �                     "@�       �                   �Z@��
ц��?             :@������������������������       �                      @�       �                   �a@      �?             8@�       �                    �?�z�G��?             $@������������������������       �                     �?�       �                   �j@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                   c@X�Cc�?             ,@������������������������       �                     @�       �                   `@X�<ݚ�?             "@������������������������       �                      @�       �                   �c@����X�?             @������������������������       �                     @�       �                    d@      �?             @������������������������       �                     �?�       �                   0d@�q�q�?             @������������������������       �                     �?�       �                    h@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   ``@�W�{�5�?B            �W@�       �                    �?����Q8�?1            �Q@�       �                   �m@���7�?.            �P@�       �                   @^@�O4R���?'            �J@�       �                   �\@Pa�	�?            �@@������������������������       �        	             &@�       �                     �?���7�?             6@������������������������       �                     @�       �                    �?�IєX�?             1@������������������������       �                     �?�       �                   pa@      �?             0@�       �                   Pi@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             ,@������������������������       �                     4@�       �                   �m@8�Z$���?             *@�       �                    d@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   0n@ףp=
�?             $@������������������������       �                     @�       �                   pn@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             8@������������������������       �                     "@�       �                   �`@��S���?             .@�       �                   �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�z�G��?             $@������������������������       �                     @�       �                    k@      �?             @�       �                   `f@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �h@ �q�q�?             8@�       �                   0g@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     (@�                          �?Ph�e���?Q            �`@�                         �_@և���X�?            �H@�                         `o@؇���X�?             5@�                           �?���Q��?             @������������������������       �                      @                        �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @                        0q@      �?             0@                        �p@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@	      
                  �p@X�Cc�?             <@������������������������       �                     @                        `a@��<b���?             7@                        �a@      �?             0@                        ``@�q�q�?             @������������������������       �                     �?                        �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@                        pd@և���X�?             @������������������������       �                      @                        �t@���Q��?             @������������������������       �                     @������������������������       �                      @      9                   @*�s���?4             U@      (                  �p@����!�?2            �T@                        pb@d��0u��?             >@                        p@�<ݚ�?             "@                         �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @       '                  �p@��s����?             5@!      "                    �?�X�<ݺ?             2@������������������������       �                     @#      $                  �p@��S�ۿ?
             .@������������������������       �                     (@%      &                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @)      0                  �a@$�q-�?             J@*      /                   �?����X�?             @+      ,                  pa@�q�q�?             @������������������������       �                     @-      .                  a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?1      8                  �^@`Ӹ����?            �F@2      7                  �q@@4և���?             <@3      6                   �?8�Z$���?             *@4      5                  `c@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �        
             .@������������������������       �                     1@������������������������       �                      @;      L                   �?�G�z��?'             N@<      E                  �s@��R[s�?            �A@=      B                   �?HP�s��?             9@>      ?                   e@�nkK�?             7@������������������������       �                     4@@      A                  `m@�q�q�?             @������������������������       �                      @������������������������       �                     �?C      D                  �b@      �?              @������������������������       �                     �?������������������������       �                     �?F      G                   �?�z�G��?             $@������������������������       �                      @H      K                   c@      �?              @I      J                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @M      ^                   �? �o_��?             9@N      Q                  �g@�GN�z�?             6@O      P                  �e@�q�q�?             @������������������������       �                     �?������������������������       �                      @R      ]                  @g@�S����?             3@S      X                  �d@�����H�?             2@T      W                  �l@@4և���?
             ,@U      V                  �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@Y      Z                  p@      �?             @������������������������       �                      @[      \                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?_      `                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMaKK�r�  hR�B        u@     �x@      4@     �_@      2@     �_@      0@     �J@      @     �B@              @      @     �@@      @      3@      @      ,@               @      @      (@      @      (@      �?      (@              @      �?      @      �?                      @       @              �?                      @      @      ,@      �?      ,@      �?                      ,@       @              "@      0@      "@      "@              @      "@      @              @      "@      @      "@      �?      @               @      �?              �?       @                       @              @       @     �R@              @       @     �P@              E@       @      9@       @      $@               @       @       @               @       @                      .@       @             �s@     �p@      R@     �d@     �A@      &@      (@      $@      @      @               @      @      @              @      @      �?       @              �?      �?      �?                      �?      "@      @       @      @      @      �?       @      �?       @                      �?      @               @       @              �?       @      �?       @                      �?      �?      �?              �?      �?              7@      �?      7@                      �?     �B@     @c@      @       @      @                       @      ?@      c@      �?      8@              (@      �?      (@              $@      �?       @               @      �?              >@      `@      &@      Z@      &@      W@              7@      &@     @Q@      $@     @Q@      @     �J@      @      ?@      �?      *@      �?      "@              @      �?      @      �?      @      �?      �?              �?      �?                      @              �?              @      @      2@      �?      0@              ,@      �?       @      �?                       @      @       @      @                       @              6@      @      0@      @      "@      @      @      �?      �?              �?      �?               @      @       @       @       @                       @              �?      �?      @      �?       @               @      �?                      @      �?      @      �?      �?      �?                      �?              @      �?                      (@      3@      8@      2@      $@      .@      $@      .@      @      @      �?      @      �?      @                      �?       @              "@      @      @      @      �?               @      @       @       @      �?              �?       @               @      �?                      @      @                      @      @              �?      ,@      �?      @      �?                      @              &@     �n@      Z@     `k@     �Q@     ``@      :@      [@      9@      8@      ,@      7@      (@      "@              ,@      (@       @              (@      (@      @      @              �?      @       @      @                       @      @      "@              @      @      @               @      @       @      @               @       @              �?       @      �?      �?              �?      �?              �?      �?              �?       @      �?                       @      U@      &@     �P@      @     �O@      @      J@      �?      @@      �?      &@              5@      �?      @              0@      �?      �?              .@      �?      �?      �?              �?      �?              ,@              4@              &@       @       @      �?              �?       @              "@      �?      @              @      �?              �?      @              @      �?      �?              @      �?      @                      �?      1@      @      "@               @      @      �?      @              @      �?              @      @      @              @      @      @      �?      @                      �?               @      7@      �?      &@      �?      &@                      �?      (@              V@     �F@      5@      <@      @      2@       @      @               @       @      �?              �?       @              �?      .@      �?      @              @      �?                      $@      2@      $@              @      2@      @      ,@       @      �?       @              �?      �?      �?      �?                      �?      *@              @      @       @               @      @              @       @             �P@      1@     �P@      .@      3@      &@       @      @       @       @       @                       @              @      1@      @      1@      �?      @              ,@      �?      (@               @      �?       @                      �?              @      H@      @      @       @      @       @      @              �?       @      �?                       @      �?             �E@       @      :@       @      &@       @      @       @      @                       @      @              .@              1@                       @      ;@     �@@      "@      :@       @      7@      �?      6@              4@      �?       @               @      �?              �?      �?              �?      �?              @      @               @      @      �?       @      �?              �?       @              @              2@      @      1@      @      �?       @      �?                       @      0@      @      0@       @      *@      �?       @      �?              �?       @              &@              @      �?       @              �?      �?      �?                      �?              �?      �?       @      �?                       @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ��fbhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfMUhgh"h#K �r�  h%�r�  Rr�  (KMU�r�  hn�B�J         t                   �`@�#i����?�           ��@       E                    �?����m�?�            �r@                            �?�r����?�             l@       	                   �`@��S���?	             .@                          @^@؇���X�?             @������������������������       �                     @                           `@�q�q�?             @������������������������       �                     �?������������������������       �                      @
                          �^@      �?              @������������������������       �                     @������������������������       �                     �?       .                    �?\�����?�            @j@                           �?�NW���?k            �c@                          �h@�FVQ&�?            �@@                          �g@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     9@       '                    �?�[|x��?T            �_@       &                   �a@h�˹�?6             S@       !                   �[@�X�C�?'             L@                          �_@      �?             0@������������������������       �                     @                          `k@      �?	             (@                          �Z@z�G�z�?             @������������������������       �                     @������������������������       �                     �?                           �`@����X�?             @                           `@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @"       #                   `_@��(\���?             D@������������������������       �                     >@$       %                   0j@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     4@(       )                   �p@p���?             I@������������������������       �                    �G@*       -                   `_@�q�q�?             @+       ,                   x{@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?/       D                    �?��[�8��?!            �I@0       ;                   �b@     ��?             @@1       :                   Pl@      �?             4@2       3                   �X@�n_Y�K�?
             *@������������������������       �                      @4       7                   �k@���!pc�?             &@5       6                    `@؇���X�?             @������������������������       �                     �?������������������������       �                     @8       9                    `@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @<       ?                   �c@      �?             (@=       >                    S@      �?             @������������������������       �                     @������������������������       �                     �?@       A                   @e@      �?              @������������������������       �                     �?B       C                   �q@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     3@F       a                   @\@�s��:��?6             S@G       N                     �?      �?             8@H       M                   `c@���Q��?             @I       J                   �m@�q�q�?             @������������������������       �                     �?K       L                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @O       `                    a@���y4F�?             3@P       [                   @Y@      �?             0@Q       V                    �?և���X�?             @R       S                    �?�q�q�?             @������������������������       �                     �?T       U                   `X@      �?              @������������������������       �                     �?������������������������       �                     �?W       Z                   �T@      �?             @X       Y                   @\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?\       ]                   �l@�����H�?             "@������������������������       �                     @^       _                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @b       q                    �?��
ц��?#             J@c       d                   �]@V������?            �B@������������������������       �                     "@e       h                     �?��>4և�?             <@f       g                    �?      �?             @������������������������       �                     @������������������������       �                     @i       n                   �c@���|���?             6@j       m                   @L@����X�?             @k       l                   P`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @o       p                    @z�G�z�?
             .@������������������������       �                     (@������������������������       �                     @r       s                   �q@�r����?             .@������������������������       �                     *@������������������������       �                      @u       �                    I@F�Q�j�?           {@v       �                   @e@r�q��?             H@w       �                    �?�ʈD��?            �E@x       y                   �U@`Jj��?             ?@������������������������       �                     �?z                          �^@(;L]n�?             >@{       ~                   Pa@$�q-�?	             *@|       }                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �        	             1@�       �                    �?r�q��?             (@������������������������       �                     �?�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                    `@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �g@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       
                  �c@x�(�3��?�            x@�       �                   pa@�4�[<��?�             j@�       �                   r@>A�F<�?             C@�       �                     �?<���D�?            �@@������������������������       �                     @�       �                    �?8�Z$���?             :@�       �                    �?���y4F�?             3@�       �                   �`@���Q��?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �`@@4և���?	             ,@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                     @�       �                    b@���Q��?             @�       �                   hs@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �l@X�<ݚ�?h            `e@�       �                   @c@�4F����?-            �T@�       �                    �?��ga�=�?&            �P@�       �                     �?�jTM��?"            �N@�       �                    �?@4և���?             ,@������������������������       �                     �?������������������������       �                     *@�       �                    �?p�v>��?            �G@�       �                    �?П[;U��?             =@�       �                   �j@8�A�0��?             6@�       �                    i@�E��ӭ�?             2@�       �                   `h@�q�q�?             (@�       �                   �b@�z�G��?             $@�       �                   �e@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   @b@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �?�X�<ݺ?             2@������������������������       �                      @�       �                   �j@ףp=
�?             $@������������������������       �                     @�       �                    b@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    _@������?             .@�       �                    g@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    b@r�q��?             (@������������������������       �                     @�       �                     �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                     �?��9܂�?;            @V@�       �                   �a@|��?���?             ;@�       �                    �?؇���X�?             @������������������������       �                     @�       �                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �r@��Q��?             4@�       �                   �p@      �?	             0@�       �                    b@      �?              @�       �                   �n@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �a@      �?             @�       �                   y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�                          a@�U���?)             O@�       �                   �r@H�z�G�?             D@�       �                   0c@��.k���?             A@�       �                    _@X�<ݚ�?             ;@�       �                   `o@�t����?             1@�       �                   �b@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?"pc�
�?             &@�       �                   �p@�<ݚ�?             "@������������������������       �                     @�       �                    ]@�q�q�?             @������������������������       �                     @�       �                   Pb@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?�z�G��?             $@�       �                   �`@���Q��?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �\@؇���X�?             @�       �                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�                           t@r�q��?             @������������������������       �                     @������������������������       �                     �?                        c@�C��2(�?             6@                        pc@P���Q�?             4@������������������������       �                     (@                        8p@      �?              @������������������������       �                     �?������������������������       �                     @      	                  r@      �?              @������������������������       �                     �?������������������������       �                     �?      N                  �r@"pc�
�?i             f@      ?                  �e@V��~��?[            �b@      >                  �r@������?A            @Z@      #                   �?j�*�'�?@            �Y@                        �d@և���X�?             <@                        `a@X�<ݚ�?
             2@                         �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @                         �?      �?              @������������������������       �                      @                         b@�q�q�?             @                         j@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @      "                  Pe@z�G�z�?             $@                          �?�����H�?             "@������������������������       �                     �?      !                   e@      �?              @                         �d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?$      )                  �\@�r����?/            �R@%      &                   �?X�<ݚ�?             "@������������������������       �                     @'      (                   �?r�q��?             @������������������������       �                     �?������������������������       �                     @*      3                   �?�C��2(�?,            �P@+      2                  �e@z�G�z�?             4@,      1                  d@�����H�?             2@-      .                  �_@�<ݚ�?             "@������������������������       �                     �?/      0                  �c@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                      @4      5                  �n@�nkK�?             G@������������������������       �                     >@6      =                  0a@      �?             0@7      <                  �p@z�G�z�?             $@8      9                  �o@�q�q�?             @������������������������       �                     �?:      ;                  �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @@      A                    �?��S�ۿ?            �F@������������������������       �                     ,@B      M                   @��a�n`�?             ?@C      L                   �?��S�ۿ?             >@D      K                   �?@4և���?             <@E      F                  0j@����X�?             @������������������������       �                     �?G      H                   �?r�q��?             @������������������������       �                     @I      J                  pf@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        
             5@������������������������       �                      @������������������������       �                     �?O      T                   �? ��WV�?             :@P      Q                  �r@؇���X�?             @������������������������       �                     @R      S                   �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             3@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMUKK�r�  hR�BP       `u@     �x@      P@     �m@      >@     `h@      @       @      @      �?      @               @      �?              �?       @              �?      @              @      �?              7@     `g@      (@     `b@       @      ?@       @      @              @       @                      9@      $@      ]@      "@     �P@      "@     �G@      @      $@              @      @      @      �?      @              @      �?              @       @       @       @       @                       @      @              @     �B@              >@      @      @      @                      @              4@      �?     �H@             �G@      �?       @      �?      �?      �?                      �?              �?      &@      D@      &@      5@      @      .@      @       @       @              @       @      �?      @      �?                      @       @       @               @       @                      @      @      @      @      �?      @                      �?      @      @              �?      @      @      @                      @              3@      A@      E@      @      2@       @      @       @      �?      �?              �?      �?              �?      �?                       @      @      .@      @      (@      @      @      �?       @              �?      �?      �?              �?      �?               @       @      �?       @      �?                       @      �?              �?       @              @      �?      �?              �?      �?                      @      <@      8@      :@      &@      "@              1@      &@      @      @      @                      @      ,@       @       @      @       @      @       @                      @               @      (@      @      (@                      @       @      *@              *@       @             `q@     `c@       @      D@      @     �C@       @      =@      �?              �?      =@      �?      (@      �?      �?      �?                      �?              &@              1@       @      $@      �?              �?      $@              @      �?      @               @      �?      �?              �?      �?              @      �?      @                      �?     �p@     �\@     �_@     �T@      ?@      @      =@      @      @              6@      @      .@      @       @      @               @       @      �?              �?       @              *@      �?      �?      �?      �?                      �?      (@              @               @      @      �?      @              @      �?              �?             �W@      S@      L@      :@      J@      .@      G@      .@      *@      �?              �?      *@             �@@      ,@      0@      *@      *@      "@      *@      @      @      @      @      @      @      �?              �?      @                       @               @      @                      @      @      @              @      @              1@      �?       @              "@      �?      @              @      �?              �?      @              @              @      &@       @      �?              �?       @               @      $@              @       @      @              @       @             �C@      I@      ,@      *@      �?      @              @      �?      �?              �?      �?              *@      @      (@      @      @      @      @      �?      @                      �?              @       @              �?      @      �?      �?      �?                      �?               @      9@     �B@      7@      1@      2@      0@      (@      .@      @      (@      @      @      @                      @       @      "@       @      @              @       @      @              @       @      �?       @                      �?               @      @      @      @       @      @      �?              �?      @                      �?      @      �?              �?      @              @      �?      �?      �?      �?                      �?      @              @      �?      @                      �?       @      4@      �?      3@              (@      �?      @      �?                      @      �?      �?      �?                      �?      b@      @@     �]@      ?@     @S@      <@     @S@      :@      (@      0@      $@       @       @       @       @                       @       @      @               @       @      @       @      �?              �?       @                      @       @       @      �?       @              �?      �?      @      �?      @              @      �?                      @      �?             @P@      $@      @      @              @      @      �?              �?      @              N@      @      0@      @      0@       @      @       @              �?      @      �?      @                      �?      "@                       @      F@       @      >@              ,@       @       @       @      �?       @              �?      �?      �?              �?      �?              @              @                       @      E@      @      ,@              <@      @      <@       @      :@       @      @       @              �?      @      �?      @               @      �?       @                      �?      5@               @                      �?      9@      �?      @      �?      @              @      �?              �?      @              3@        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ$�phG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r   (hKhfMhgh"h#K �r  h%�r  Rr  (KM�r  hn�B=         &                   �_@"��G,�?�           ��@                           �?��˥W1�?V            `a@                           �?��.��?%            �N@                          `]@@4և���?             <@������������������������       �                     *@                          @b@�r����?
             .@                          �`@$�q-�?             *@                           I@z�G�z�?             @	       
                   �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                          �c@      �?              @������������������������       �                     �?������������������������       �                     �?                            �?r٣����?            �@@������������������������       �                     �?                           \@     ��?             @@������������������������       �                      @                           �?�q�q�?             8@������������������������       �                     @                          �`@�KM�]�?             3@������������������������       �                     ,@                          @]@���Q��?             @������������������������       �                      @������������������������       �                     @                           �? ���J��?1            �S@������������������������       �        !             I@       %                   p`@@4և���?             <@                             �?�r����?	             .@������������������������       �                     �?!       "                    `@؇���X�?             ,@������������������������       �                      @#       $                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     *@'       �                    �?@�����?h           ��@(       �                   �b@��N�[�?�             s@)       �                   0f@$��fF?�?�            @o@*       +                   �Q@0u��A��?�             n@������������������������       �                      @,       1                   @Z@��&�F"�?�            �m@-       0                    �?�q�q�?             @.       /                   `l@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @2       I                     �?>���Rp�?�             m@3       8                   `_@p�ݯ��?             C@4       7                    Z@$�q-�?             *@5       6                   �l@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@9       >                    �?�q�����?             9@:       =                    b@�q�q�?             "@;       <                   y@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @?       D                   @m@      �?	             0@@       C                    k@r�q��?             @A       B                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @E       H                    �?ףp=
�?             $@F       G                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @J       K                   `d@v�9�z��?q            @h@������������������������       �                     �?L       a                    _@���[�A�?p             h@M       T                   `l@ �Cc}�?/             U@N       O                   pk@��Y��]�?            �D@������������������������       �                     =@P       Q                    �?�8��8��?             (@������������������������       �                     "@R       S                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @U       V                   �l@&^�)b�?            �E@������������������������       �                     @W       X                    Z@��-�=��?            �C@������������������������       �                     0@Y       Z                    �?�㙢�c�?             7@������������������������       �                     @[       `                    `@���y4F�?             3@\       ]                   �Z@�q�q�?             @������������������������       �                      @^       _                   �[@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        	             *@b       q                   0i@"��3؞�?A            @[@c       n                   �`@X�<ݚ�?
             2@d       m                   �h@�	j*D�?             *@e       f                    f@ףp=
�?             $@������������������������       �                     @g       h                    �?r�q��?             @������������������������       �                     @i       l                    g@�q�q�?             @j       k                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @o       p                   �f@z�G�z�?             @������������������������       �                     �?������������������������       �                     @r       �                   �b@8�Z$���?7            �V@s       t                   �k@�����H�?1            @T@������������������������       �                     5@u       �                    �?R���Q�?%             N@v       w                    �?�:pΈ��?             I@������������������������       �        
             0@x       y                   0l@H�V�e��?             A@������������������������       �                     �?z       {                    a@"pc�
�?            �@@������������������������       �                     $@|                          �n@��+7��?             7@}       ~                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @_@z�G�z�?	             4@������������������������       �                     &@�       �                   pd@X�<ݚ�?             "@�       �                   �p@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   ``@z�G�z�?             $@������������������������       �                     @�       �                   pq@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?      �?             $@�       �                   �n@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     $@�       �                   @^@@3����?             K@�       �                    f@ 7���B�?             ;@������������������������       �                     8@�       �                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ;@�       �                   �_@�q4���?�            0r@�       �                   pn@F�����?             �L@�       �                   @]@X�Cc�?             E@�       �                    �?���B���?             :@�       �                   @_@�IєX�?	             1@�       �                   @\@؇���X�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                   @a@X�<ݚ�?             "@������������������������       �                      @�       �                    [@����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?      �?             0@�       �                   �c@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       �                   `^@������?
             .@�       �                   �p@���|���?             &@������������������������       �                     @�       �                   �\@և���X�?             @�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �l@:�&���?�            @m@�       �                   d@������?>            @V@�       �                     �?և���X�?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     �?�       �                    b@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                     �?������?9            �T@������������������������       �                     8@�       �                    �? 	��p�?&             M@������������������������       �                     ;@�       �                    �?��� ��?             ?@�       �                   a@ �Cc}�?             <@�       �                   �j@�nkK�?             7@������������������������       �        	             1@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �d@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       
                   �?>���Rp�?[             b@�       �                   pm@d}h���?N            �_@�       �                    @�q�q�?             (@�       �                    �?X�<ݚ�?             "@������������������������       �                      @�       �                   �b@և���X�?             @������������������������       �                     @�       �                   �l@      �?             @������������������������       �                      @�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    ]@r�q��?F            �\@�       �                     �?�eP*L��?             &@������������������������       �                     @�       �                   0n@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                     �?�`�=	�??            �Y@�       �                   0a@`Ql�R�?            �G@������������������������       �                     ;@�       �                   0r@P���Q�?             4@�       �                    @؇���X�?             @�       �                    b@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@�       	                   f@4և����?$             L@�                          d@�rF���?#            �K@�       �                   b@^������?            �A@�       �                    �?�����H�?	             2@�       �                   �o@z�G�z�?             $@������������������������       �                     @�       �                   �p@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   0o@j���� �?             1@�       �                   �m@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �b@�	j*D�?             *@������������������������       �                     @                         �c@      �?              @                         �?z�G�z�?             @                        c@      �?             @                         b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@������������������������       �                     �?                        �o@D�n�3�?             3@                        0o@�����H�?             "@                        �n@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                          �?�z�G��?             $@������������������������       �                     �?                         �?�<ݚ�?             "@                        �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @r  tr  bh�h"h#K �r  h%�r  Rr	  (KMKK�r
  hR�Bp       @s@     �z@      (@     �_@      $@     �I@       @      :@              *@       @      *@      �?      (@      �?      @      �?      @              @      �?                      �?               @      �?      �?      �?                      �?       @      9@      �?              @      9@               @      @      1@      @               @      1@              ,@       @      @       @                      @       @      S@              I@       @      :@       @      *@              �?       @      (@               @       @      @              @       @                      *@     �r@     �r@     @R@     �l@      R@     @f@      O@     @f@       @              N@     @f@      @       @      �?       @      �?                       @      @              L@      f@      8@      ,@      (@      �?      @      �?              �?      @              "@              (@      *@      @      @      @      �?      @                      �?               @      @      $@      @      �?      �?      �?              �?      �?              @              �?      "@      �?      @              @      �?                       @      @@     @d@      �?              ?@     @d@      "@     �R@      �?      D@              =@      �?      &@              "@      �?       @      �?                       @       @     �A@      @              @     �A@              0@      @      3@              @      @      .@      @       @       @               @       @               @       @                      *@      6@     �U@       @      $@      @      "@      �?      "@              @      �?      @              @      �?       @      �?      �?              �?      �?                      �?      @              @      �?              �?      @              ,@     @S@      "@      R@              5@      "@     �I@      @     �E@              0@      @      ;@      �?              @      ;@              $@      @      1@       @      �?       @                      �?      @      0@              &@      @      @      @      @              @      @                       @       @       @              @       @       @       @                       @      @      @      @       @               @      @                      @      $@              �?     �J@      �?      :@              8@      �?       @      �?                       @              ;@     �k@      Q@      ?@      :@      ;@      .@      5@      @      0@      �?      @      �?      @              �?      �?      �?                      �?      $@              @      @               @      @       @               @      @              @      $@      @      �?              �?      @                      "@      @      &@      @      @              @      @      @      �?      @              @      �?              @                      @      h@      E@     �T@      @      @      @      �?              @      @      �?               @      @              @       @             �S@      @      8@              K@      @      ;@              ;@      @      9@      @      6@      �?      1@              @      �?      @                      �?      @       @               @      @               @      �?              �?       @             �[@     �A@     �X@      ;@      @       @      @      @               @      @      @      @              �?      @               @      �?      �?              �?      �?                      @     �W@      3@      @      @      @              �?      @      �?                      @     @V@      ,@      G@      �?      ;@              3@      �?      @      �?      @      �?      �?      �?      �?                      �?       @              @              *@             �E@      *@     �E@      (@      7@      (@      0@       @       @       @      @              @       @               @      @               @              @      $@      @      �?              �?      @              @      "@              @      @      @      @      �?      @      �?      �?      �?      �?                      �?       @              �?                      @      4@                      �?      &@       @       @      �?      @      �?      @                      �?      @              @      @      �?               @      @       @      �?       @                      �?              @r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJW:+LhG        hNhG        h8Kh9Kh:h"h#K �r  h%�r  Rr  (KK�r  hR�C              �?r  tr  bhFhVhAC       r  �r  Rr  hZKh[h\Kh"h#K �r  h%�r  Rr  (KK�r  hA�C       r  tr  bK�r  Rr  }r   (hKhfMhgh"h#K �r!  h%�r"  Rr#  (KM�r$  hn�B�=         �                    �?�#i����?�           ��@                          �c@�^����?�            �w@       
                   P`@`�q�0ܴ?E            �W@                          �b@�k~X��?6             R@������������������������       �        .            �O@       	                   �c@�����H�?             "@                           S@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?��2(&�?             6@                           �?և���X�?             @������������������������       �                     �?                            �?      �?             @������������������������       �                     �?                          `b@���Q��?             @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        
             .@       U                   n@PQr,���?�            �q@       N                   �a@v�`����?Q            @^@       =                   ``@�Pf����?A            �W@       :                   �m@�E����?0             R@       9                   d@
��[��?,            @P@                           @X@d��0u��?'             N@                          @_@����X�?             @                          �l@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?!       "                   Pf@f1r��g�?$            �J@������������������������       �                     $@#       4                    �?&^�)b�?            �E@$       '                    g@z�G�z�?             >@%       &                   @_@      �?             @������������������������       �                     �?������������������������       �                     @(       -                    `@ȵHPS!�?             :@)       ,                   `i@�IєX�?             1@*       +                   �h@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             (@.       /                   �j@�<ݚ�?             "@������������������������       �                     �?0       1                    _@      �?              @������������������������       �                     @2       3                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?5       6                   �l@8�Z$���?             *@������������������������       �                     "@7       8                   �\@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @;       <                    �?����X�?             @������������������������       �                      @������������������������       �                     @>       M                   �c@8����?             7@?       L                   0c@b�2�tk�?             2@@       I                    �?ҳ�wY;�?             1@A       B                   �i@�θ�?             *@������������������������       �                     @C       D                   �Y@      �?             @������������������������       �                      @E       H                   @_@      �?             @F       G                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @J       K                   �j@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @O       P                    �?$�q-�?             :@������������������������       �                      @Q       R                   �`@�����H�?             2@������������������������       �                     (@S       T                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     @V       k                    a@ޭ�W[��?a            @d@W       j                   �`@�ʈD��?4            �U@X       _                   �p@4�2%ޑ�?            �A@Y       Z                   �[@X�<ݚ�?             "@������������������������       �                     @[       \                    �?�q�q�?             @������������������������       �                     �?]       ^                   `o@���Q��?             @������������������������       �                      @������������������������       �                     @`       a                    U@8�Z$���?             :@������������������������       �                     �?b       e                    �?H%u��?             9@c       d                     �?�}�+r��?             3@������������������������       �                     �?������������������������       �        
             2@f       i                     �?�q�q�?             @g       h                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                    �I@l       �                   �a@\�Uo��?-             S@m       z                     �?\�����?            �K@n       u                   �r@���|���?             6@o       p                   `b@r�q��?             (@������������������������       �                     @q       t                   @o@����X�?             @r       s                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @v       y                    �?���Q��?             $@w       x                   0c@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @{       �                    `@���|���?            �@@|       �                    f@z�G�z�?             4@}       �                   �^@�����H�?
             2@~                           ]@"pc�
�?             &@������������������������       �                     @�       �                   �p@�q�q�?             @������������������������       �                      @�       �                   Pb@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   `a@�n_Y�K�?             *@�       �                   ``@�z�G��?             $@�       �                   �q@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   Xt@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �d@��s����?             5@�       �                    �?�X�<ݺ?             2@������������������������       �                      @�       �                    f@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @�       �                   �c@t�F�}�?�            Pv@�       �                    `@�X���?             F@�       �                    �?؇���X�?             ,@������������������������       �                      @�       �                     �?r�q��?
             (@������������������������       �                     �?�       �                    `@�C��2(�?	             &@������������������������       �                     @�       �                    \@r�q��?             @�       �                   �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   `@*;L]n�?             >@������������������������       �        	             *@�       �                    �?������?	             1@�       �                   �a@����X�?             ,@������������������������       �                      @�       �                   pb@�q�q�?             @������������������������       �                      @�       �                   �d@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?��k�0��?�            �s@�       �                   @\@��%F��?V             a@�       �                    Z@���Q��?             $@�       �                    X@z�G�z�?             @������������������������       �                      @�       �                   `Y@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    [@���Q��?             @������������������������       �                      @�       �                     �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   d@4Jı@�?P            �_@�       �                     �?$�Z����?0             S@������������������������       �                     =@�       �                   p@��|�5��?            �G@�       �                    �?      �?             @@������������������������       �                     8@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �                   �q@�q�q�?             .@�       �                   �c@�eP*L��?	             &@�       �                    �?      �?              @�       �                   Xp@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �I@�       �                     �?v�X��?k             f@�       �                   `X@PN��T'�?!             K@�       �                   �k@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �? i���t�?            �H@������������������������       �                     4@�       �                    �?д>��C�?             =@�       �                   �`@�J�4�?             9@������������������������       �        
             *@�       �                   a@�q�q�?             (@������������������������       �                      @������������������������       �                     @�       �                   @_@      �?             @������������������������       �                      @�       �                   `]@      �?              @������������������������       �                     �?������������������������       �                     �?�                          @�-ῃ�?J            �^@�                          �?2E�=<��?=            �X@�       �                   �`@JyK���?4            �U@�       �                    ]@X�;�^o�?             �K@�       �                   `\@      �?
             4@�       �                   �[@r�q��?	             2@�       �                    �?�8��8��?             (@������������������������       �                     �?�       �                   @[@�C��2(�?             &@�       �                   @Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    `@ >�֕�?            �A@�       �                   �g@ףp=
�?             4@������������������������       �                     �?�       �                   `k@�}�+r��?
             3@�       �                   �i@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@������������������������       �                     .@�                          �f@      �?             @@�       �                   0d@"pc�
�?             &@�       �                    d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                        �d@�q�q�?             5@                        pc@��S�ۿ?	             .@������������������������       �                     &@                        �c@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                         �?�eP*L��?	             &@	                        �n@և���X�?             @
                        P`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                        0b@      �?             @������������������������       �                     @������������������������       �                     �?                         o@      �?             8@                        �j@�	j*D�?             *@������������������������       �                     @                         �?      �?              @                         �?      �?             @������������������������       �                     �?������������������������       �                     @                         �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@r%  tr&  bh�h"h#K �r'  h%�r(  Rr)  (KMKK�r*  hR�B�       `u@     �x@     �T@     `r@      @     �V@      �?     �Q@             �O@      �?       @      �?      �?      �?                      �?              @      @      3@      @      @              �?      @      @              �?      @       @      �?       @      �?                       @       @                      .@     �S@     �i@     �D@      T@     �C@      L@      7@     �H@      2@     �G@      *@     �G@      @       @      @       @      @                       @      �?               @     �F@              $@       @     �A@      @      8@      @      �?              �?      @              @      7@      �?      0@      �?      @              @      �?                      (@       @      @      �?              �?      @              @      �?       @               @      �?               @      &@              "@       @       @       @                       @      @              @       @               @      @              0@      @      &@      @      &@      @      $@      @      @              @      @       @              �?      @      �?      �?              �?      �?                       @      �?      @              @      �?                      �?      @               @      8@               @       @      0@              (@       @      @       @                      @      C@      _@       @     �S@       @      ;@      @      @              @      @       @      �?              @       @               @      @              @      6@      �?              @      6@      �?      2@      �?                      2@       @      @       @       @       @                       @               @             �I@      >@      G@      :@      =@      ,@       @      $@       @      @              @       @      �?       @               @      �?              @              @      @      @      @              @      @                       @      (@      5@      @      0@       @      0@       @      "@              @       @      @               @       @       @       @                       @              @       @               @      @      @      @      @      @              @      @               @              �?       @               @      �?              @      1@      �?      1@               @      �?      "@              "@      �?              @             0p@     �X@      .@      =@       @      (@               @       @      $@      �?              �?      $@              @      �?      @      �?       @               @      �?                      @      *@      1@              *@      *@      @      $@      @       @               @      @               @       @       @       @                       @      @             �n@     @Q@      ^@      1@      @      @      �?      @               @      �?       @      �?                       @      @       @       @              �?       @               @      �?              ]@      &@     @P@      &@      =@              B@      &@      ?@      �?      8@              @      �?      @                      �?      @      $@      @      @      @      @      @      @              @      @              �?                      @              @     �I@              _@      J@      G@       @       @      @       @                      @      F@      @      4@              8@      @      5@      @      *@               @      @       @                      @      @      �?       @              �?      �?              �?      �?             �S@      F@     @Q@      =@      P@      7@      H@      @      .@      @      .@      @      &@      �?      �?              $@      �?      �?      �?      �?                      �?      "@              @       @               @      @                       @     �@@       @      2@       @              �?      2@      �?      @      �?      @                      �?      .@              .@              0@      0@      "@       @      �?       @               @      �?               @              @      ,@      �?      ,@              &@      �?      @      �?                      @      @              @      @      @      @      �?      @              @      �?              @              �?      @              @      �?              "@      .@      "@      @      @              @      @      �?      @      �?                      @      @      �?      @                      �?              &@r+  tr,  bubhhubh)�r-  }r.  (hhh	h
hNhKhKhG        hh hNhJF<KdhG        hNhG        h8Kh9Kh:h"h#K �r/  h%�r0  Rr1  (KK�r2  hR�C              �?r3  tr4  bhFhVhAC       r5  �r6  Rr7  hZKh[h\Kh"h#K �r8  h%�r9  Rr:  (KK�r;  hA�C       r<  tr=  bK�r>  Rr?  }r@  (hKhfMOhgh"h#K �rA  h%�rB  RrC  (KMO�rD  hn�BHI         (                   @E@�#i����?�           ��@                           �?��|,��?L             _@                           �?����"$�?8            �U@                           �?XB���?'             M@                          @^@�����H�?             2@������������������������       �                      @������������������������       �                     0@������������������������       �                     D@	                          �b@�>4և��?             <@
                          `[@P���Q�?             4@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@                           �?      �?              @������������������������       �                     @������������������������       �                     @                          @\@p�ݯ��?             C@������������������������       �                     @                           �?     ��?             @@������������������������       �                     @       '                    @l��[B��?             =@                           �?��
ц��?             :@                           �?և���X�?             @������������������������       �                     �?                           �?      �?             @������������������������       �                     @������������������������       �                     @       &                   pb@�\��N��?	             3@       %                    `@�θ�?             *@       "                    �?և���X�?             @        !                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @#       $                   �]@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @)       �                   �a@��t��?�           �@*       q                   �`@6�Vp�?           �|@+       .                   �V@�����C�?h             d@,       -                    q@r�q��?             @������������������������       �                     @������������������������       �                     �?/       F                     �?���]�?e            `c@0       =                    �?V������?            �B@1       4                    �?�J�4�?             9@2       3                   �`@      �?              @������������������������       �                     @������������������������       �                     @5       6                    �?�IєX�?             1@������������������������       �                      @7       8                    �?�����H�?             "@������������������������       �                     �?9       <                   �q@      �?              @:       ;                   �l@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @>       E                   �s@�q�q�?             (@?       D                   �`@      �?              @@       C                    �?      �?             @A       B                   @_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @G       H                   �X@F�4�Dj�?N            �]@������������������������       �        
             2@I       J                   @Y@H.�!���?D             Y@������������������������       �                     @K       l                    �?L� P?)�?A            @X@L       c                    �?`K�����?3            @R@M       ^                    �?�X�C�?'             L@N       ]                   �p@ i���t�?"            �H@O       \                   �`@؇���X�?            �A@P       Q                    �?      �?             @@������������������������       �                     .@R       [                   `o@�t����?             1@S       T                   `_@      �?             0@������������������������       �                     &@U       V                   @Y@z�G�z�?             @������������������������       �                     �?W       Z                   �k@      �?             @X       Y                    `@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@_       b                    k@և���X�?             @`       a                   �g@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @d       k                   P`@��.k���?             1@e       j                   �\@�	j*D�?	             *@f       i                    @և���X�?             @g       h                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @m       n                   pa@ �q�q�?             8@������������������������       �                     2@o       p                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?r       �                   �l@�����?�            �r@s       �                    �?j��>��?S            ``@t       u                     �?�ʻ����?             A@������������������������       �                     @v       {                   Pe@      �?             >@w       z                   @`@؇���X�?             @x       y                   �_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @|       �                   ``@�û��|�?             7@}       �                    g@"pc�
�?             &@~                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    a@�q�q�?             (@������������������������       �                     @�       �                   �h@r�q��?             @�       �                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �`@DE�SA_�?>            @X@�       �                   �a@ �q�q�?.             R@�       �                   Pg@z�G�z�?
             .@������������������������       �                     @�       �                   Pa@�z�G��?             $@������������������������       �                     @�       �                    �?      �?             @�       �                   �g@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �        $            �L@�       �                    �?z�G�z�?             9@�       �                    @�GN�z�?             6@�       �                   �c@�����H�?             2@�       �                   @b@����X�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                    a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   0m@X���Og�?d            �d@�       �                     �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                   hq@�X����?]            @c@�       �                    �?T��?:            �Y@�       �                   Pa@���@M^�?             ?@������������������������       �                     @�       �                   ``@l��
I��?             ;@�       �                   �n@      �?             0@������������������������       �                     �?�       �                   �a@��S���?
             .@������������������������       �                      @�       �                   @[@��
ц��?	             *@������������������������       �                      @�       �                    �?���|���?             &@�       �                     �?և���X�?             @������������������������       �                     @�       �                   �^@      �?             @�       �                    \@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   @_@      �?             @�       �                   @p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                     �?O�o9%�?)            �Q@������������������������       �                     .@�       �                    c@4և����?             L@�       �                    �?�q�q�?             8@�       �                    _@�G�z��?             4@�       �                   �\@z�G�z�?             $@������������������������       �                     @�       �                   �p@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    a@ףp=
�?             $@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �o@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �p@     ��?             @@������������������������       �                     ;@�       �                    @���Q��?             @�       �                    �?�q�q�?             @�       �                   Pd@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                     �?��
ц��?#             J@�       �                   @b@r�q��?
             (@������������������������       �                      @������������������������       �                     $@�       �                    �?�G�z��?             D@�       �                   pe@�Gi����?            �B@�       �                   @[@r�q��?             8@������������������������       �                     �?�       �                   �_@�LQ�1	�?             7@������������������������       �                     (@�       �                   pa@���!pc�?             &@�       �                   �`@�q�q�?             @�       �                   xs@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     @�       �                   @c@z�G�z�?             @�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?8�Z$���?             *@�       �                    f@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     @�       <                   �?ҳ�wY;�?e             c@�       �                   `e@*;L]n�?Q             ^@�       �                    �?����X�?             @������������������������       �                      @������������������������       �                     @�                           �?�d�
t��?L            @\@�                          �?X�<ݚ�?             B@�                         �w@*;L]n�?             >@�                         �s@��}*_��?             ;@                          �?\X��t�?             7@                        @a@z�G�z�?             $@                        �^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @                        �c@8�Z$���?             *@                         �?����X�?             @������������������������       �                      @	                         @���Q��?             @
                        �g@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @                         �?      �?             @������������������������       �                     @������������������������       �                     @                        �a@����X�?6            @S@                         �?և���X�?             @������������������������       �                      @                          @���Q��?             @                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                        �b@��R[s�?2            �Q@������������������������       �        
             *@      3                  �n@�����?(            �L@      *                   �?�g�y��?             ?@       '                  0l@      �?             0@!      &                   k@@4և���?	             ,@"      %                   �?؇���X�?             @#      $                  `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @(      )                   �?      �?              @������������������������       �                     �?������������������������       �                     �?+      2                  �b@�r����?             .@,      1                   c@      �?              @-      .                  �`@�q�q�?             @������������������������       �                     �?/      0                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @4      7                  �p@ȵHPS!�?             :@5      6                  xp@      �?              @������������������������       �                     @������������������������       �                      @8      9                  �r@�X�<ݺ?             2@������������������������       �                     &@:      ;                   �?؇���X�?             @������������������������       �                     @������������������������       �                     �?=      H                   �?�'�`d�?            �@@>      E                  �e@�KM�]�?             3@?      D                   �?�IєX�?
             1@@      A                  �r@�8��8��?             (@������������������������       �                     $@B      C                  �w@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @F      G                  �q@      �?              @������������������������       �                     �?������������������������       �                     �?I      N                  �a@X�Cc�?             ,@J      M                   �?ףp=
�?             $@K      L                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @rE  trF  bh�h"h#K �rG  h%�rH  RrI  (KMOKK�rJ  hR�B�       `u@     �x@      5@     �Y@      @     �S@       @      L@       @      0@       @                      0@              D@      @      7@      �?      3@      �?      �?      �?                      �?              2@      @      @      @                      @      ,@      8@              @      ,@      2@              @      ,@      .@      ,@      (@      @      @      �?              @      @      @                      @      $@      "@      $@      @      @      @      �?       @      �?                       @      @      �?              �?      @              @                      @              @     t@     r@     �p@     �g@     �J@      [@      @      �?      @                      �?      H@     �Z@      :@      &@      5@      @      @      @      @                      @      0@      �?       @               @      �?      �?              @      �?      @      �?      @                      �?      @              @      @      @      @      @      @      @      �?      @                      �?               @       @                      @      6@      X@              2@      6@     �S@      @              3@     �S@      2@     �K@      "@     �G@      @      F@      @      >@       @      >@              .@       @      .@      �?      .@              &@      �?      @              �?      �?      @      �?      �?      �?                      �?               @      �?              @                      ,@      @      @      @      �?              �?      @                       @      "@       @      "@      @      @      @      @      �?              �?      @                      @      @                      @      �?      7@              2@      �?      @              @      �?             �j@     �T@      [@      7@      3@      .@      @              .@      .@      @      �?      @      �?      @                      �?       @              "@      ,@       @      "@       @      �?              �?       @                       @      @      @      @              �?      @      �?      �?      �?                      �?              @     @V@       @     @Q@      @      (@      @      @              @      @      @              �?      @      �?       @               @      �?                      �?     �L@              4@      @      1@      @      0@       @      @       @      @              �?       @      �?                       @      &@              �?      @              @      �?              @             �Z@     �M@      �?      $@      �?                      $@     @Z@     �H@     @S@      9@      3@      (@              @      3@       @       @       @      �?              @       @               @      @      @               @      @      @      @      @      @              �?      @      �?      �?              �?      �?                       @      @      �?      �?      �?      �?                      �?       @              &@              M@      *@      .@             �E@      *@      ,@      $@      &@      "@       @       @              @       @      @              @       @              "@      �?      @               @      �?              �?       @              @      �?      @                      �?      =@      @      ;@               @      @       @      �?      �?      �?              �?      �?              �?                       @      <@      8@      $@       @               @      $@              2@      6@      .@      6@      @      4@      �?              @      4@              (@      @       @       @      �?      �?      �?              �?      �?              �?              �?      @              @      �?      @      �?      �?      �?                      �?              @      &@       @      �?       @               @      �?              $@              @              K@     �X@     �G@     @R@      @       @               @      @              E@     �Q@      4@      0@      1@      *@      1@      $@      *@      $@       @       @       @       @               @       @                      @      &@       @      @       @       @              @       @      �?       @               @      �?               @              @              @                      @      @      @              @      @              6@     �K@      @      @       @               @      @       @      �?              �?       @                       @      2@      J@              *@      2@     �C@      .@      0@       @      ,@      �?      *@      �?      @      �?       @      �?                       @              @              @      �?      �?      �?                      �?      *@       @      @       @      �?       @              �?      �?      �?              �?      �?              @              @              @      7@       @      @              @       @              �?      1@              &@      �?      @              @      �?              @      :@       @      1@      �?      0@      �?      &@              $@      �?      �?      �?                      �?              @      �?      �?      �?                      �?      @      "@      �?      "@      �?      �?      �?                      �?               @      @        rK  trL  bubhhubh)�rM  }rN  (hhh	h
hNhKhKhG        hh hNhJؽ�hG        hNhG        h8Kh9Kh:h"h#K �rO  h%�rP  RrQ  (KK�rR  hR�C              �?rS  trT  bhFhVhAC       rU  �rV  RrW  hZKh[h\Kh"h#K �rX  h%�rY  RrZ  (KK�r[  hA�C       r\  tr]  bK�r^  Rr_  }r`  (hKhfM?hgh"h#K �ra  h%�rb  Rrc  (KM?�rd  hn�B�E         �                   �`@�/�$�y�?�           ��@       s                    �?R�����?�            @v@                            �?��7;k�?�            Pp@                          �v@�	j*D�?             J@                          @e@�GN�z�?             F@       	                   �Z@RB)��.�?            �E@                          �r@      �?              @������������������������       �                     @������������������������       �                     @
                           _@(N:!���?            �A@������������������������       �                     ,@                           �?��s����?             5@                          @]@      �?             @������������������������       �                     �?                           `@���Q��?             @������������������������       �                     �?                          �_@      �?             @                          `^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           ^@��S�ۿ?             .@������������������������       �                     "@                          �^@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                          �z@      �?              @������������������������       �                     @������������������������       �                      @       V                    �?f�D;��?�             j@        K                   P`@�����H�?`             c@!       2                    �?����1�?Y            @b@"       1                   �k@�f�¦ζ?A            �Z@#       (                    \@h�WH��?#             K@$       %                    �?�q�q�?             @������������������������       �                     �?&       '                   �h@      �?              @������������������������       �                     �?������������������������       �                     �?)       .                    `@�IєX�?             �I@*       -                   �Y@`Ql�R�?            �G@+       ,                   �X@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                    �C@/       0                   @`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                    �J@3       <                   �_@�θ�?            �C@4       ;                    ]@�q�q�?             "@5       :                   �^@؇���X�?             @6       7                    \@      �?             @������������������������       �                      @8       9                   @V@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @=       B                    S@ףp=
�?             >@>       ?                   `]@z�G�z�?             $@������������������������       �                     @@       A                    ^@�q�q�?             @������������������������       �                      @������������������������       �                     �?C       D                   �p@P���Q�?             4@������������������������       �                     *@E       F                   �]@؇���X�?             @������������������������       �                      @G       H                   �e@z�G�z�?             @������������������������       �                      @I       J                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @L       M                   p`@և���X�?             @������������������������       �                     �?N       O                   �`@�q�q�?             @������������������������       �                      @P       Q                   �Z@      �?             @������������������������       �                     �?R       S                   �`@�q�q�?             @������������������������       �                     �?T       U                    b@      �?              @������������������������       �                     �?������������������������       �                     �?W       X                   @\@>4և���?!             L@������������������������       �                     @Y       `                    \@䯦s#�?            �J@Z       [                   �_@�����?	             5@������������������������       �                     ,@\       _                    �?����X�?             @]       ^                   Pi@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @a       b                   P`@     ��?             @@������������������������       �                     @c       d                   @]@� �	��?             9@������������������������       �                     @e       h                    �?�z�G��?             4@f       g                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?i       r                    @������?             1@j       k                   �a@      �?
             0@������������������������       �                     "@l       q                    _@և���X�?             @m       p                   �^@      �?             @n       o                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?t       �                   Xr@�:nR&y�??            �W@u       v                    f@h�����?7             U@������������������������       �                     F@w       x                     �?��(\���?             D@������������������������       �                     �?y       �                    �?�7��?            �C@z       {                    ^@�����?             5@������������������������       �        
             *@|       }                    �?      �?              @������������������������       �                     �?~                          �k@����X�?             @������������������������       �                     @�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     2@�       �                   @^@���|���?             &@������������������������       �                     @������������������������       �                     @�                          �?������?�            �w@�       �                   �c@6P��[�?�            �t@�       �                   �g@ާb�y��?r            �g@�       �                   Pa@">�֕�?            �A@������������������������       �                     @�       �                   Pd@      �?             @@�       �                    @���Q��?	             .@�       �                   @E@      �?             (@�       �                     �?���Q��?             $@������������������������       �                     @�       �                   c@և���X�?             @�       �                    d@�q�q�?             @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �b@�t����?	             1@�       �                   �e@      �?              @������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@�       �                   8q@���Q��?^            `c@�       �                     �?�e�,��?E            �]@�       �                   �a@`Jj��?             ?@������������������������       �                     0@�       �                    �?�r����?	             .@�       �                   po@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �                    �?�f7�z�?4            �U@�       �                    �?4�2%ޑ�?            �A@�       �                   �b@      �?              @�       �                    c@r�q��?             @�       �                   pb@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �i@�+$�jP�?             ;@������������������������       �                     �?�       �                    �?8�Z$���?             :@�       �                   �j@��S�ۿ?             .@�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@�       �                   Pm@���!pc�?             &@������������������������       �                      @������������������������       �                     @�       �                    c@D>�Q�?              J@�       �                    �?���!pc�?            �@@�       �                   `o@z�G�z�?             4@������������������������       �                     *@�       �                   �_@և���X�?             @������������������������       �                     @�       �                   �`@      �?             @������������������������       �                      @�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �a@�n_Y�K�?             *@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �                    @���Q��?             @�       �                   �b@      �?             @������������������������       �                     �?�       �                   0m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@�       �                   �b@^H���+�?            �B@�       �                   0a@r�q��?             8@�       �                    a@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�����?             5@������������������������       �                     .@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                     �?z�G�z�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                     �?�	j*D�?             *@������������������������       �                      @�       �                    c@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�                         q@�7��ެ�?Y            `a@�       �                     �?,�T�6�?A             Z@������������������������       �                     C@�       �                   �d@r�q��?-            �P@�       �                    o@�X����?             6@�       �                    ]@      �?             4@������������������������       �                     @�       �                    �?�t����?             1@������������������������       �                     "@�       �                    �?      �?              @������������������������       �                     @�       �                   Pd@�q�q�?             @������������������������       �                     �?�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�                         �b@�C��2(�?             F@�                         �f@@4և���?             E@�                          @�C��2(�?            �@@�                         �`@ 	��p�?             =@�                         ``@�t����?             1@�                          �?      �?             0@�                          0k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             *@������������������������       �                     �?������������������������       �                     (@                        0f@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@	      
                  �c@      �?              @������������������������       �                     �?������������������������       �                     �?                          �?^������?            �A@                        s@����X�?             @                         �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                        �_@X�Cc�?             <@                        pe@      �?	             (@                         �?�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @                        �r@      �?
             0@                         �?z�G�z�?             @������������������������       �                     @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@                         �Z@���Q �?&            �H@������������������������       �                     @!      "                  0a@�D����?"             E@������������������������       �                     @#      *                   �?4�B��?            �B@$      )                   n@և���X�?             @%      &                   `@      �?             @������������������������       �                      @'      (                  �g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @+      0                   �?�z�G��?             >@,      -                  ``@�IєX�?             1@������������������������       �                     $@.      /                  Pa@؇���X�?             @������������������������       �                     �?������������������������       �                     @1      2                  `b@�n_Y�K�?             *@������������������������       �                     �?3      4                   _@�q�q�?
             (@������������������������       �                     @5      6                  �O@      �?              @������������������������       �                     �?7      >                   �?և���X�?             @8      ;                    �?      �?             @9      :                  @q@�q�q�?             @������������������������       �                      @������������������������       �                     �?<      =                  �e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?re  trf  bh�h"h#K �rg  h%�rh  Rri  (KM?KK�rj  hR�B�        t@     �y@     �T@     q@      S@      g@      B@      0@      A@      $@      A@      "@      @      @              @      @              ?@      @      ,@              1@      @      @      @              �?      @       @              �?      @      �?      �?      �?      �?                      �?       @              ,@      �?      "@              @      �?              �?      @                      �?       @      @              @       @              D@      e@      1@      a@      ,@     �`@      @     �Y@      @     �H@       @      �?      �?              �?      �?              �?      �?              @      H@      �?      G@      �?      @              @      �?                     �C@       @       @               @       @                     �J@      "@      >@      @      @      @      �?      @      �?       @              �?      �?      �?                      �?      @                       @      @      ;@       @       @              @       @      �?       @                      �?      �?      3@              *@      �?      @               @      �?      @               @      �?       @      �?                       @      @      @      �?               @      @               @       @       @              �?       @      �?      �?              �?      �?              �?      �?              7@     �@@      @              4@     �@@       @      3@              ,@       @      @       @      @       @                      @               @      2@      ,@      @              &@      ,@      @              @      ,@       @      �?       @                      �?      @      *@      @      (@              "@      @      @      �?      @      �?      �?              �?      �?                       @      @                      �?      @      V@      @     @T@              F@      @     �B@      �?               @     �B@       @      3@              *@       @      @              �?       @      @              @       @      �?       @                      �?              2@      @      @      @                      @     �m@     �a@     �k@     @[@      Z@     �U@      &@      8@      @               @      8@      @      "@      @      @      @      @              @      @      @      @       @       @       @               @       @               @                      �?       @                      @       @      .@       @      @              @       @       @       @                       @              "@     @W@      O@      T@      C@      =@       @      0@              *@       @      @       @               @      @              "@             �I@      B@       @      ;@      @      @      �?      @      �?       @               @      �?                      @       @              @      6@      �?              @      6@      �?      ,@      �?       @      �?                       @              (@      @       @               @      @             �E@      "@      8@      "@      0@      @      *@              @      @              @      @      �?       @              �?      �?              �?      �?               @      @      @              @      @              @      @       @      @      �?      �?               @      �?       @                      �?              �?      3@              *@      8@      @      4@       @      �?              �?       @               @      3@              .@       @      @      �?              �?      @      �?       @      �?                       @               @      "@      @       @              �?      @      �?                      @      ]@      7@     @W@      &@      C@             �K@      &@      .@      @      .@      @              @      .@       @      "@              @       @      @              �?       @              �?      �?      �?      �?                      �?               @      D@      @     �C@      @      >@      @      ;@       @      .@       @      .@      �?       @      �?              �?       @              *@                      �?      (@              @      �?              �?      @              "@              �?      �?              �?      �?              7@      (@      @       @      �?       @               @      �?              @              2@      $@      @      @      @      @              @      @              @              (@      @      �?      @              @      �?      �?              �?      �?              &@              1@      @@              @      1@      9@      @              (@      9@      @      @      @      �?       @              �?      �?              �?      �?                      @      "@      5@      �?      0@              $@      �?      @      �?                      @       @      @              �?       @      @      @              @      @              �?      @      @      @      @      �?       @               @      �?               @      �?       @                      �?      �?        rk  trl  bubhhubh)�rm  }rn  (hhh	h
hNhKhKhG        hh hNhJX��vhG        hNhG        h8Kh9Kh:h"h#K �ro  h%�rp  Rrq  (KK�rr  hR�C              �?rs  trt  bhFhVhAC       ru  �rv  Rrw  hZKh[h\Kh"h#K �rx  h%�ry  Rrz  (KK�r{  hA�C       r|  tr}  bK�r~  Rr  }r�  (hKhfMhgh"h#K �r�  h%�r�  Rr�  (KM�r�  hn�B=         �                    �?���
%�?�           ��@       �                   �y@b�h�d.�?�            x@       |                    �?v�}��?�            �w@       E                   `a@��G�<�?�            �q@       ,                    a@      �?h             e@                           �?�"�q��?7            �W@       
                   0i@���7�?             6@       	                   �g@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             .@                          �[@��oh���?(            @R@                            �?�G��l��?             5@                           Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?X�<ݚ�?             2@                           [@��
ц��?	             *@                          �_@���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @                          �Z@���Q��?             @������������������������       �                      @                          �Y@�q�q�?             @������������������������       �                     �?������������������������       �                      @       !                     �?ȵHPS!�?             J@                          �_@      �?             @������������������������       �                     �?                            i@�q�q�?             @������������������������       �                     �?������������������������       �                      @"       #                   �]@�8��8��?             H@������������������������       �                     2@$       +                    I@�r����?             >@%       (                    �?���|���?             &@&       '                   `]@؇���X�?             @������������������������       �                     @������������������������       �                     �?)       *                   P`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             3@-       >                    �?F��}��?1            @R@.       7                   �c@`'�J�?"            �I@/       6                   �[@�(\����?             D@0       5                   �a@�}�+r��?             3@1       2                     �?؇���X�?             @������������������������       �                     @3       4                   �Z@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@������������������������       �                     5@8       =                   �d@�C��2(�?             &@9       <                    o@؇���X�?             @:       ;                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @?       D                    S@�C��2(�?             6@@       A                   `]@�q�q�?             @������������������������       �                     @B       C                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     0@F       W                     �?.��$�?D            @]@G       N                   pn@��Zy�?            �C@H       M                   e@X�Cc�?
             ,@I       J                    �?r�q��?             @������������������������       �                     �?K       L                   `T@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @O       V                   0d@`�Q��?             9@P       Q                    `@��s����?	             5@������������������������       �                     @R       U                   �`@�X�<ݺ?             2@S       T                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     .@������������������������       �                     @X       {                   �f@R�}e�.�?/            �S@Y       Z                   �Z@�+e�X�?-            �R@������������������������       �                      @[       x                   pc@��oh���?+            @R@\       ]                    �?�#ʆA��?            �J@������������������������       �                     $@^       w                   0c@8�$�>�?            �E@_       p                    �?�(�Tw��?            �C@`       g                   pj@     ��?             @@a       b                   �a@���Q��?             $@������������������������       �                     @c       d                   @b@z�G�z�?             @������������������������       �                     @e       f                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?h       m                   r@��2(&�?             6@i       j                   �a@      �?	             0@������������������������       �                     (@k       l                   @b@      �?             @������������������������       �                     �?������������������������       �                     @n       o                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     @q       v                   `b@����X�?             @r       s                   Pm@r�q��?             @������������������������       �                     @t       u                   �n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @y       z                   �t@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?������������������������       �                     @}       �                   @s@��8�$>�?D            @X@~       �                    �?�==Q�P�?B            �W@       �                   �^@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@�       �                   �l@ ��N8�?;             U@������������������������       �        /            �P@�       �                   �\@�X�<ݺ?             2@�       �                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             0@�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    `@Z�L[IZ�?�            �u@�       �                   P`@d��0u��?:            �V@�       �                    a@hP�vCu�?            �D@�       �                    \@�r����?             .@������������������������       �                     @�       �                    �?�<ݚ�?             "@�       �                   @^@      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �?ȵHPS!�?             :@�       �                    �?HP�s��?             9@�       �                    Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   xt@�X�<ݺ?             2@������������������������       �        
             1@������������������������       �                     �?������������������������       �                     �?�       �                   c@ZՏ�m|�?!            �H@�       �                   @]@      �?             0@�       �                   �W@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             ,@�       �                     �?�'�`d�?            �@@������������������������       �                     @�       �                    g@ܷ��?��?             =@�       �                   pd@@4և���?             <@������������������������       �                     �?�       �                   �p@ 7���B�?             ;@������������������������       �                     5@�       �                   �a@r�q��?             @������������������������       �                     @�       �                    q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                     �?�����=�?�            0p@�       �                   �Q@0�>���?:            �V@������������������������       �                      @�       �                   �`@X;��?9            @V@������������������������       �        )            �P@�       �                   �`@��2(&�?             6@�       �                    �?���Q��?             @������������������������       �                      @�       �                   @q@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   `c@�IєX�?             1@������������������������       �        	             *@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?\`*�s�?k             e@�       �                   pq@h�˹�?.             S@�       �                   @a@���U�?#            �L@�       �                   �a@@�E�x�?            �H@�       �                   @_@@4և���?	             ,@�       �                   (p@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@������������������������       �                    �A@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �                    b@p�ݯ��?             3@�       �                    _@�C��2(�?             &@�       �                    d@      �?              @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?      �?              @�       �                    �?���Q��?             @������������������������       �                     �?�       �                   `c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   `a@�+Fi��?=             W@������������������������       �        	             ,@�       �                   �b@a��t��?4            �S@�       �                   �a@��<b���?             7@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?R���Q�?	             4@������������������������       �                     @�       �                   �`@d}h���?             ,@�       �                   0m@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @�                         Pp@�b��[��?)            �K@�                         �d@���X�K�?            �F@�       �                   �f@�n_Y�K�?             :@������������������������       �                     @�                          �?      �?             4@�       �                   @Y@      �?
             0@������������������������       �                      @�                          b@����X�?	             ,@�       �                    �?�θ�?             *@�       �                    @�q�q�?             @�       �                   pn@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   @^@؇���X�?             @������������������������       �                      @�                          �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        `e@�S����?             3@������������������������       �                     @                         f@      �?
             (@                        �`@�q�q�?             @      	                   �?�q�q�?             @������������������������       �                     �?
                         _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        `]@r�q��?             @������������������������       �                     �?������������������������       �                     @                        pf@���Q��?
             $@                         \@      �?              @������������������������       �                     �?                        0c@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hR�Bp       0s@     �z@     �P@     �s@     �O@     �s@     �M@     @l@      5@     `b@      1@     �S@      �?      5@      �?      @              @      �?                      .@      0@     �L@      $@      &@       @      �?              �?       @               @      $@      @      @      @      @              @      @                      @       @      @               @       @      �?              �?       @              @      G@       @       @      �?              �?       @      �?                       @      @      F@              2@      @      :@      @      @      �?      @              @      �?              @      �?      @                      �?              3@      @     @Q@       @     �H@      �?     �C@      �?      2@      �?      @              @      �?      @              @      �?                      (@              5@      �?      $@      �?      @      �?      �?      �?                      �?              @              @       @      4@       @      @              @       @      �?              �?       @                      0@      C@     �S@      1@      6@      "@      @      �?      @              �?      �?      @              @      �?               @               @      1@      @      1@      @              �?      1@      �?       @               @      �?                      .@      @              5@     �L@      2@     �L@       @              0@     �L@      .@      C@              $@      .@      <@      &@      <@      "@      7@      @      @      @              �?      @              @      �?      �?      �?                      �?      @      3@      �?      .@              (@      �?      @      �?                      @       @      @       @                      @       @      @      �?      @              @      �?      �?      �?                      �?      �?              @              �?      3@              3@      �?              @              @     @W@      @      W@       @      "@       @                      "@      �?     �T@             �P@      �?      1@      �?      �?              �?      �?                      0@      �?      �?              �?      �?              @              n@      [@     �@@     �L@      9@      0@       @      *@              @       @      @       @      @       @      �?              �?       @                      @              �?      7@      @      7@       @      @      �?              �?      @              1@      �?      1@                      �?              �?       @     �D@      �?      .@      �?      �?              �?      �?                      ,@      @      :@      @              @      :@       @      :@      �?              �?      :@              5@      �?      @              @      �?       @      �?                       @      �?              j@     �I@     �U@      @               @     �U@      @     �P@              3@      @      @       @       @              �?       @               @      �?              0@      �?      *@              @      �?      @                      �?     �^@      G@     �P@      "@     �K@       @      H@      �?      *@      �?      @      �?      @                      �?      $@             �A@              @      �?      @                      �?      (@      @      $@      �?      @      �?      �?      �?      �?                      �?      @              @               @      @       @      @              �?       @       @               @       @                      @     �K@     �B@      ,@             �D@     �B@      @      2@       @      �?       @                      �?      @      1@              @      @      &@      @      @      @                      @               @      B@      3@      @@      *@      0@      $@      @              $@      $@      @      $@       @              @      $@      @      $@       @      @      �?      @              @      �?              �?              �?      @               @      �?      @              @      �?              �?              @              0@      @      @              "@      @      @       @      �?       @              �?      �?      �?      �?                      �?      @              @      �?              �?      @              @      @       @      @      �?              �?      @      �?                      @       @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ���EhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfMAhgh"h#K �r�  h%�r�  Rr�  (KMA�r�  hn�B8F                            �?�r,��?�           ��@       �                    �?�;n���?x           X�@       @                   P`@¦	^_�?�            `s@       	                     �?Z�J�p�?h            �d@                          �`@j���� �?             1@������������������������       �                     "@                          �_@      �?              @������������������������       �                     @������������������������       �                     �?
                           �?(E����?]            �b@                          �a@��FM ò?B            @Z@                          �`@�IєX�?/             Q@                          `_@`���i��?             F@������������������������       �                     B@                          �\@      �?              @                          �k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                          �e@      �?             8@������������������������       �                     "@                          �Y@z�G�z�?	             .@������������������������       �                      @                          i@$�q-�?             *@������������������������       �                     �?������������������������       �                     (@������������������������       �                    �B@       '                   �_@�zv�X�?             F@                          �X@������?             .@������������������������       �                     �?                            [@d}h���?             ,@������������������������       �                     @!       &                   �Z@      �?              @"       %                   �q@      �?             @#       $                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @(       ;                    _@V�a�� �?             =@)       ,                    X@�J�4�?             9@*       +                   @V@�q�q�?             @������������������������       �                      @������������������������       �                     �?-       2                    S@��2(&�?             6@.       /                   `]@�<ݚ�?             "@������������������������       �                     @0       1                   �]@      �?             @������������������������       �                      @������������������������       �                      @3       4                   �]@$�q-�?             *@������������������������       �                     @5       :                   @^@؇���X�?             @6       7                   �c@r�q��?             @������������������������       �                     @8       9                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?<       ?                   �b@      �?             @=       >                    `@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?A       �                   `f@�a�2���?U             b@B       u                   �b@h+�v:�?O             a@C       t                   pb@X3_��?+            �Q@D       M                     �?�ՙ/�?(            �O@E       F                   �]@���Q��?             $@������������������������       �                     @G       H                   �X@؇���X�?             @������������������������       �                     @I       L                    c@      �?             @J       K                   a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?N       a                   �^@䯦s#�?#            �J@O       Z                   �]@p�ݯ��?             3@P       Q                    a@�q�q�?             "@������������������������       �                     �?R       S                   �W@      �?              @������������������������       �                     �?T       U                    �?����X�?             @������������������������       �                      @V       Y                   �\@���Q��?             @W       X                   �n@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?[       \                   a@ףp=
�?             $@������������������������       �                     �?]       ^                   Pk@�����H�?             "@������������������������       �                     @_       `                   �p@      �?             @������������������������       �                     �?������������������������       �                     @b       i                   �f@������?             A@c       d                   �`@�q�q�?             "@������������������������       �                     �?e       h                    U@      �?              @f       g                   `b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @j       q                    �?HP�s��?             9@k       l                    �?���N8�?             5@������������������������       �                     @m       n                    b@��S�ۿ?
             .@������������������������       �                     (@o       p                   �e@�q�q�?             @������������������������       �                     �?������������������������       �                      @r       s                   r@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @v       �                    �?�	j*D�?$            @P@w       z                   �n@"pc�
�?             6@x       y                    _@      �?             @������������������������       �                     �?������������������������       �                     @{       |                   �u@�X�<ݺ?
             2@������������������������       �                     *@}       ~                    a@z�G�z�?             @������������������������       �                     @       �                   pc@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �\@�lg����?            �E@������������������������       �                     ,@�       �                     �?П[;U��?             =@�       �                    a@�<ݚ�?             "@������������������������       �                     @�       �                   @e@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?�G�z��?             4@�       �                    d@j���� �?             1@������������������������       �                     @�       �                   �k@��
ц��?             *@������������������������       �                     @�       �                   �_@�z�G��?             $@������������������������       �                      @�       �                    b@      �?              @�       �                   0a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @b@      �?              @������������������������       �                     @������������������������       �                     �?�                         c@��%W��?�            Pq@�       �                    �?�/g�+�?�            @o@�       �                    �?�u��R�?H            �Z@�       �                     �?D�n�3�?             3@������������������������       �                     @�       �                   �m@�q�q�?             (@������������������������       �                     @�       �                   �r@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    �?����!p�?<             V@�       �                    I@��S�ۿ?4            �R@�       �                   `_@      �?             @������������������������       �                      @������������������������       �                      @�       �                   e@0z�(>��?1            �Q@�       �                   l@=QcG��?!            �G@������������������������       �                     4@�       �                   0m@�����H�?             ;@������������������������       �                     �?�       �                    b@$�q-�?             :@�       �                   �^@���N8�?             5@�       �                     �?ףp=
�?             $@������������������������       �                     @�       �                   �c@؇���X�?             @������������������������       �                     @�       �                    d@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                   �a@z�G�z�?             @������������������������       �                      @�       �                   @q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     8@������������������������       �                     *@�       �                   P`@�f|��?_            �a@�       �                    �?.p����??            @Y@�       �                   �[@H��?"�?4             U@�       �                    a@p�ݯ��?             3@�       �                   `^@؇���X�?             @������������������������       �                     @�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �X@�8��8��?	             (@������������������������       �                     �?������������������������       �                     &@�       �                     �?����?'            @P@������������������������       �                     ;@�       �                   �m@�KM�]�?             C@�       �                   �m@�㙢�c�?             7@�       �                   �g@��2(&�?             6@�       �                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�KM�]�?             3@�       �                   �]@      �?             @������������������������       �                      @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    ^@��S�ۿ?	             .@������������������������       �                     �?������������������������       �                     ,@������������������������       �                     �?������������������������       �        	             .@�       �                   �c@j���� �?             1@�       �                   @j@�q�q�?             (@�       �                   �\@����X�?             @������������������������       �                     �?�       �                    @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �a@և���X�?              E@�       �                   �`@և���X�?             <@������������������������       �                     @�       �                   �d@      �?             8@�       �                   pi@�t����?             1@�       �                    �?����X�?             @������������������������       �                     �?�       �                    �?r�q��?             @�       �                    T@�q�q�?             @������������������������       �                     �?�       �                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     @�                          �b@؇���X�?
             ,@�       �                   pb@����X�?             @�       �                   `_@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @      	                    �?�5��?             ;@                        Pg@      �?             $@������������������������       �                     @                        @e@����X�?             @������������������������       �                     @                        �u@�q�q�?             @������������������������       �                     �?������������������������       �                      @
                        pc@ҳ�wY;�?             1@������������������������       �                     �?                        �`@     ��?             0@                        �l@և���X�?             @                         �?      �?             @������������������������       �                     �?                        �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                        @g@�����H�?             "@������������������������       �                      @������������������������       �                     �?      6                  �a@��
CJ�?X            `b@      %                   �?�uw\l��?7            @W@                        ``@�i�y�?%            �O@������������������������       �                    �G@      "                   �?      �?             0@                        �^@$�q-�?             *@������������������������       �                     "@                        0a@      �?             @������������������������       �                      @       !                  @a@      �?              @������������������������       �                     �?������������������������       �                     �?#      $                   `@�q�q�?             @������������������������       �                      @������������������������       �                     �?&      5                   @���Q��?             >@'      .                  �`@����"�?             =@(      -                  pa@r�q��?             (@)      ,                   �?�C��2(�?             &@*      +                  �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?/      0                  �m@�IєX�?
             1@������������������������       �                     &@1      2                  �`@r�q��?             @������������������������       �                     @3      4                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?7      8                  Pc@ 7���B�?!             K@������������������������       �                     4@9      :                  �b@�IєX�?             A@������������������������       �                     *@;      <                  �e@�����?             5@������������������������       �                     �?=      >                  �^@P���Q�?             4@������������������������       �                     &@?      @                   a@�����H�?             "@������������������������       �                     �?������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMAKK�r�  hR�B       �t@     Py@     0s@     �q@     �V@     �k@      ?@     �`@      $@      @      "@              �?      @              @      �?              5@      `@      @     @Y@      @      P@      �?     �E@              B@      �?      @      �?       @      �?                       @              @      @      5@              "@      @      (@       @              �?      (@      �?                      (@             �B@      1@      ;@      &@      @              �?      &@      @      @              @      @      �?      @      �?      �?              �?      �?                       @      @              @      7@      @      5@      �?       @               @      �?              @      3@       @      @              @       @       @       @                       @      �?      (@              @      �?      @      �?      @              @      �?      �?      �?                      �?              �?       @       @       @      �?       @                      �?              �?     �M@     @U@      J@      U@      @@     �C@      8@     �C@      @      @      @              �?      @              @      �?      @      �?       @      �?                       @              �?      4@     �@@      (@      @      @      @              �?      @      @      �?               @      @               @       @      @       @       @       @                       @              �?      "@      �?      �?               @      �?      @              @      �?              �?      @               @      :@      @      @              �?      @       @       @       @               @       @              @               @      7@      �?      4@              @      �?      ,@              (@      �?       @      �?                       @      �?      @              @      �?               @              4@     �F@      @      2@      @      �?              �?      @              �?      1@              *@      �?      @              @      �?      �?              �?      �?              0@      ;@              ,@      0@      *@      @       @      @              �?       @               @      �?              "@      &@      @      $@              @      @      @              @      @      @               @      @      �?      @      �?      @                      �?      @               @      �?              �?       @              @      �?      @                      �?      k@      N@      i@     �H@     �W@      *@      &@       @      @              @       @      @              �?       @               @      �?             �T@      @     �Q@      @       @       @               @       @              Q@      @      F@      @      4@              8@      @              �?      8@       @      4@      �?      "@      �?      @              @      �?      @              @      �?              �?      @              &@              @      �?       @               @      �?       @                      �?      8@              *@             �Z@      B@     �T@      2@     @R@      &@      (@      @      �?      @              @      �?       @      �?                       @      &@      �?              �?      &@             �N@      @      ;@              A@      @      3@      @      3@      @       @      �?              �?       @              1@       @      @      �?       @              �?      �?              �?      �?              ,@      �?              �?      ,@                      �?      .@              $@      @      @      @      @       @              �?      @      �?      @                      �?              @      @              8@      2@      (@      0@              @      (@      (@      @      (@      @       @              �?      @      �?       @      �?      �?              �?      �?              �?      �?              @                      $@      @              (@       @      @       @      �?      �?              �?      �?              @      �?      @                      �?      @              0@      &@      @      @              @      @       @      @              �?       @      �?                       @      &@      @              �?      &@      @      @      @      @      �?      �?               @      �?              �?       @                      @       @      �?       @                      �?      6@     @_@      4@     @R@       @     �N@             �G@       @      ,@      �?      (@              "@      �?      @               @      �?      �?              �?      �?              �?       @               @      �?              2@      (@      2@      &@       @      $@      �?      $@      �?      �?      �?                      �?              "@      �?              0@      �?      &@              @      �?      @              �?      �?      �?                      �?              �?       @      J@              4@       @      @@              *@       @      3@      �?              �?      3@              &@      �?       @      �?                       @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ:9)bhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfM)hgh"h#K �r�  h%�r�  Rr�  (KM)�r�  hn�B�@         @                     �?T8���?�           ��@       3                   �c@�<ݚ��?_             b@       "                   �a@�
�G�?9             V@                           �?     ��?'             P@                           �?L紂P�?             �I@       	                   �[@������?            �D@                           c@�q�q�?             @������������������������       �                      @������������������������       �                     �?
                          @_@�˹�m��?             C@������������������������       �        	             &@                          �r@�����H�?             ;@                          �`@`2U0*��?             9@������������������������       �        
             4@                          @_@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                          �b@�z�G��?             $@������������������������       �                     @������������������������       �                     @       !                    b@�n_Y�K�?             *@                          a@      �?             $@                          �q@      �?             @������������������������       �                      @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           @�q�q�?             @������������������������       �                     @                           �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @#       ,                   �b@�q�q�?             8@$       +                   �m@@�0�!��?             1@%       &                    �?�z�G��?             $@������������������������       �                     @'       *                    `@      �?             @(       )                    X@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @-       .                    c@և���X�?             @������������������������       �                     @/       2                   �v@      �?             @0       1                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @4       9                   @[@h�����?&             L@5       8                    �?z�G�z�?             @6       7                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @:       ?                   d@���J��?!            �I@;       <                   Pp@      �?	             0@������������������������       �                      @=       >                   �q@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                    �A@A       �                    �?2� J��?p           p�@B       M                    �?h~��M�?�            �t@C       D                   �i@ 7���B�?"             K@������������������������       �                     3@E       F                   �Z@ >�֕�?            �A@������������������������       �                     �?G       L                   hp@г�wY;�?             A@H       I                   0a@��S�ۿ?             .@������������������������       �                     *@J       K                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@N       �                    �?a0�f��?�             q@O       �                   �a@z�G�z�?�             i@P       u                   @a@�!��Jh�?`            @b@Q       l                    �?n�6�Է�?O            �^@R       i                   �p@�����?5            �U@S       h                   �d@���}D�?)            �P@T       [                   p`@     ��?'             P@U       V                   �_@���H��?             E@������������������������       �                     4@W       Z                   `[@�GN�z�?             6@X       Y                   �X@      �?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     (@\       g                   Pb@���|���?             6@]       b                   @j@�q�q�?
             (@^       a                    a@؇���X�?             @_       `                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @c       d                   Pm@���Q��?             @������������������������       �                      @e       f                   @^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     @j       k                   �e@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?m       n                   �Q@�X�<ݺ?             B@������������������������       �                     �?o       t                   @[@��?^�k�?            �A@p       q                   a@      �?              @������������������������       �                     @r       s                    ]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ;@v       w                   �Z@
;&����?             7@������������������������       �                     @x       y                   �[@���Q��?             4@������������������������       �                      @z       �                   �m@X�<ݚ�?             2@{       |                   @_@��
ц��?	             *@������������������������       �                      @}       �                    i@�eP*L��?             &@~                          `c@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   e@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �a@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�>����?$             K@�       �                    d@@4և���?             E@������������������������       �                    �B@�       �                   `m@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �q@�8��8��?
             (@������������������������       �                     $@�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?������?4            �R@�       �                   �[@�㙢�c�?              G@�       �                   �p@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   pk@���H��?             E@�       �                    S@ �q�q�?             8@�       �                   `b@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     .@�       �                   �_@�<ݚ�?             2@�       �                    _@�r����?             .@�       �                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             (@�       �                    b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     <@�       (                  �g@�E�-���?�            `p@�       �                    `@�4��?�            @p@�       �                    �?�z�G��?&            �Q@�       �                   �S@�G�z��?             4@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?����X�?
             ,@�       �                   �[@z�G�z�?             $@������������������������       �                      @�       �                   �]@      �?              @�       �                   �p@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   pa@      �?             @������������������������       �                     �?�       �                   �o@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?z�G�z�?             I@�       �                    \@���|���?             &@������������������������       �                     @�       �                    @      �?              @�       �                   �Y@�q�q�?             @������������������������       �                      @�       �                   0a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                   `b@8�Z$���?            �C@�       �                   �Q@�FVQ&�?            �@@�       �                    �?�<ݚ�?             "@�       �                   @`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   @_@      �?             @�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     8@�       �                    n@�q�q�?             @������������������������       �                     @������������������������       �                      @�                         �c@Xf�?s��?o            �g@�       �                   @o@V������?=            �[@�       �                    �?b�h�d.�?'            �Q@�       �                   �`@     ��?$             P@�       �                   Pc@�����H�?            �F@�       �                    T@�ʈD��?            �E@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?�}�+r��?             C@�       �                   �m@      �?             @@�       �                   pa@h�����?             <@�       �                   Pi@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     9@�       �                   �m@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �P@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   Pd@p�ݯ��?
             3@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   @a@������?             .@������������������������       �                     @�       �                    �?���Q��?             $@������������������������       �                     @�       �                   �b@�q�q�?             @������������������������       �                     @�       �                   `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�                          @�p ��?            �D@�                         c@����e��?            �@@�       
                   �?f���M�?             ?@�       	                   �?�ՙ/�?             5@�                         �p@��Q��?             4@�       �                    �?      �?              @������������������������       �                     @                         `a@      �?             @������������������������       �                      @������������������������       �                      @                         �?�8��8��?             (@������������������������       �                     @                         �?r�q��?             @������������������������       �                     @                        �s@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?                         �?�z�G��?             $@������������������������       �                     @                        Pb@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                      @      #                   �?l{��b��?2            �S@                        pd@ >�֕�?-            �Q@                        Pd@�r����?	             .@                        �j@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@                        �j@      �?             @������������������������       �                     @������������������������       �                     �?      "                  �`@h㱪��?$            �K@                         �?      �?             @@                        ``@(;L]n�?             >@������������������������       �                     =@������������������������       �                     �?       !                   _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@$      '                   `@�<ݚ�?             "@%      &                  @e@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM)KK�r�  hR�B�       �t@     @y@     @\@      ?@     �M@      =@      J@      (@      F@      @     �B@      @       @      �?       @                      �?     �A@      @      &@              8@      @      8@      �?      4@              @      �?              �?      @                       @      @      @      @                      @       @      @      @      @      @      �?       @              �?      �?      �?                      �?       @      @              @       @      �?       @                      �?      @              @      1@      @      ,@      @      @              @      @      @      @      �?              �?      @                       @              @      @      @      @              �?      @      �?      �?      �?                      �?               @      K@       @      @      �?      �?      �?              �?      �?              @              I@      �?      .@      �?       @              @      �?              �?      @             �A@              k@     Pw@     �F@     �q@       @      J@              3@       @     �@@      �?              �?     �@@      �?      ,@              *@      �?      �?      �?                      �?              3@     �E@     �l@     �A@     �d@      ?@     �\@      3@      Z@      1@     �Q@      0@     �I@      *@     �I@      @     �B@              4@      @      1@      @      @              @      @                      (@       @      ,@       @      @      @      �?      �?      �?      �?                      �?      @               @      @               @       @      �?       @                      �?              $@      @              �?      3@              3@      �?               @      A@      �?              �?      A@      �?      @              @      �?      �?              �?      �?                      ;@      (@      &@              @      (@       @       @              $@       @      @      @               @      @      @      @      �?      @                      �?      �?      @              @      �?              @      �?              �?      @              @      I@      @     �C@             �B@      @       @               @      @              �?      &@              $@      �?      �?              �?      �?               @     �P@       @      C@      @      �?      @                      �?      @     �B@      �?      7@      �?       @               @      �?                      .@      @      ,@       @      *@       @      �?              �?       @                      (@       @      �?       @                      �?              <@     �e@     �V@     �e@      V@      5@     �H@      &@      "@      �?      @              @      �?              $@      @       @       @       @              @       @      @      �?      @                      �?              �?       @       @              �?       @      �?       @                      �?      $@      D@      @      @              @      @      @      @       @       @               @       @               @       @                       @      @     �@@       @      ?@       @      @      �?      @              @      �?              �?      @      �?      �?              �?      �?                       @              8@      @       @      @                       @     �b@     �C@     �S@     �@@      M@      (@      J@      (@      D@      @     �C@      @      @       @      @                       @      B@       @      >@       @      ;@      �?       @      �?              �?       @              9@              @      �?              �?      @              @              �?      �?              �?      �?              (@      @      �?      @      �?                      @      &@      @      @              @      @      @               @      @              @       @      �?              �?       @              @              4@      5@      4@      *@      4@      &@      *@       @      *@      @       @      @              @       @       @       @                       @      &@      �?      @              @      �?      @               @      �?       @                      �?              �?      @      @      @              @      @              @      @                       @               @     @R@      @     �P@      @      *@       @      $@      �?              �?      $@              @      �?      @                      �?     �J@       @      >@       @      =@      �?      =@                      �?      �?      �?      �?                      �?      7@              @       @      �?       @      �?                       @      @                       @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�BHzhG        hNhG        h8Kh9Kh:h"h#K �r�  h%�r�  Rr�  (KK�r�  hR�C              �?r�  tr�  bhFhVhAC       r�  �r�  Rr�  hZKh[h\Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hA�C       r�  tr�  bK�r�  Rr�  }r�  (hKhfMhgh"h#K �r�  h%�r�  Rr�  (KM�r�  hn�Bx=         n                   P`@�[��N�?�           ��@       9                    �?.5�/E-�?�            pt@       0                    �?���؅��?�            �m@                          �Z@��(�#H�?g            �d@������������������������       �                     @                           �?����8�?e            �d@������������������������       �                     @@       !                   `_@�禺f��?U            �`@	                          �Z@4�0_���?I            @\@
                          �i@p���?             I@������������������������       �                     :@                           �? �q�q�?             8@������������������������       �                     4@                          Pl@      �?             @������������������������       �                     �?������������������������       �                     @                           `@�? Da�?-            �O@                          �^@ҳ�wY;�?             1@                            �?8�Z$���?             *@������������������������       �                      @������������������������       �        	             &@������������������������       �                     @                            �?�nkK�?             G@                          �p@r�q��?             @������������������������       �                     @                          `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          `l@�(\����?             D@������������������������       �                     7@                           �l@�IєX�?             1@������������������������       �                     �?������������������������       �        
             0@"       #                   �\@�\��N��?             3@������������������������       �                      @$       %                    `@��.k���?             1@������������������������       �                     @&       +                   �j@և���X�?             ,@'       (                   `@      �?              @������������������������       �                     @)       *                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?,       /                    `@r�q��?             @-       .                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @1       8                    �?@	tbA@�?/            @Q@2       3                   ``@�(\����?             D@������������������������       �                     8@4       5                     �?      �?             0@������������������������       �                     �?6       7                    w@��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                     =@:       c                    �?*u�$��?6            �V@;       \                   `c@�9mf��?(            �O@<       [                   pb@�E��
��?"             J@=       Z                    �?(옄��?             G@>       Q                   P`@�K��&�?            �E@?       @                    a@8^s]e�?             =@������������������������       �                     @A       B                    ]@z�G�z�?             9@������������������������       �                     @C       H                    �?�d�����?             3@D       G                    �?����X�?             @E       F                    \@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @I       J                   �X@      �?             (@������������������������       �                      @K       P                   �l@ףp=
�?             $@L       M                   @Y@      �?             @������������������������       �                      @N       O                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @R       Y                    @X�Cc�?             ,@S       T                   �`@�q�q�?             (@������������������������       �                     @U       V                    �?����X�?             @������������������������       �                     �?W       X                    \@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @]       b                   �o@���!pc�?             &@^       a                    �?      �?             @_       `                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @d       i                     �? �Cc}�?             <@e       f                    [@����X�?             @������������������������       �                     @g       h                   �]@      �?             @������������������������       �                      @������������������������       �                      @j       m                    �?���N8�?             5@k       l                    d@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     (@o                         �e@؀�:M�?�            py@p       }                    I@z���ȋ�?�            `x@q       v                    �?r֛w���?             ?@r       u                    �?      �?              @s       t                   `b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @w       x                    �?�nkK�?             7@������������������������       �                     2@y       z                    ^@z�G�z�?             @������������������������       �                     @{       |                    �?      �?              @������������������������       �                     �?������������������������       �                     �?~       �                     �?��i�\>�?�            pv@       �                   �c@L紂P�?=            �Y@�       �                   �a@�<ݚ�?!             K@�       �                    �?��2(&�?             F@�       �                   �r@��-�=��?            �C@������������������������       �                     ;@�       �                    a@�q�q�?             (@�       �                   (s@�q�q�?             @������������������������       �                     @�       �                   y@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �^@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?���Q��?             $@�       �                   �t@X�<ݚ�?             "@�       �                    �?r�q��?             @������������������������       �                     @�       �                   @c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �`@ �q�q�?             H@������������������������       �                     C@�       �                   �e@z�G�z�?             $@�       �                    n@�q�q�?             @������������������������       �                      @�       �                   8q@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?`�J�4��?�            p@�       �                   8v@��%3�?>            @Y@�       �                    g@���|�?;            @X@�       �                   @_@�q�q�?             (@������������������������       �                     @������������������������       �                      @�       �                   n@z�G�z�?5            @U@�       �                   �c@�t����?            �I@�       �                    �?�������?             F@�       �                   �b@�C��2(�?            �@@�       �                   @[@�LQ�1	�?             7@������������������������       �                      @�       �                    �?���N8�?             5@������������������������       �                      @�       �                    b@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                     $@�       �                   `a@�eP*L��?             &@������������������������       �                     @�       �                   �a@      �?              @�       �                   @_@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                   �\@؇���X�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   0f@�IєX�?             A@�       �                    �?Pa�	�?            �@@�       �                   �a@      �?             @@�       �                   �p@�C��2(�?             &@������������������������       �                     @�       �                   @_@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     5@������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   @[@x�����?a            �c@�       �                   0n@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �l@��x_F-�?_             c@�       �                   �`@`-�I�w�?/             S@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�X�<ݺ?,             R@�       �                    @ 	��p�?$             M@�       �                   �k@`'�J�?             �I@�       �                    �?��<b�ƥ?             G@������������������������       �                     1@�       �                   �`@XB���?             =@������������������������       �                     ,@�       �                   0c@��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   0f@����X�?             @������������������������       �                     �?�       �                    a@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@�                          �?����?0            @S@�                          @����O��?,            �Q@�                         e@��$�4��?%            �M@�       �                    `@���j��?             G@�       �                   �a@�\��N��?             3@������������������������       �                      @�       �                    �?j���� �?             1@������������������������       �                     @�       �                   �p@�θ�?	             *@�       �                   �l@      �?             @������������������������       �                     �?�       �                   0m@���Q��?             @������������������������       �                      @�       �                    �?�q�q�?             @�       �                   �o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�                          �c@PN��T'�?             ;@�       �                    b@ȵHPS!�?             :@������������������������       �                     $@�       �                   `a@     ��?
             0@������������������������       �                      @�       �                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �        
             *@                         �?�q�q�?             (@                        �`@؇���X�?             @                         p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @	      
                   c@���Q��?             @������������������������       �                     @������������������������       �                      @                        0q@�q�q�?             @                        Pa@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                         �?������?
             1@                        @g@X�<ݚ�?             "@                         q@�q�q�?             @                         _@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hR�B�       �s@     Pz@      N@     �p@      7@     �j@      6@      b@      @              3@      b@              @@      3@     @\@      "@      Z@      �?     �H@              :@      �?      7@              4@      �?      @      �?                      @       @     �K@      @      &@       @      &@       @                      &@      @               @      F@      �?      @              @      �?       @      �?                       @      �?     �C@              7@      �?      0@      �?                      0@      $@      "@       @               @      "@              @       @      @      @      �?      @              �?      �?              �?      �?              �?      @      �?       @      �?                       @              @      �?      Q@      �?     �C@              8@      �?      .@              �?      �?      ,@              ,@      �?                      =@     �B@      K@      A@      =@      ?@      5@      9@      5@      9@      2@      4@      "@              @      4@      @      @              ,@      @      @       @      �?       @               @      �?              @              "@      @               @      "@      �?      @      �?       @              �?      �?      �?                      �?      @              @      "@      @      @              @      @       @      �?              @       @               @      @                       @              @      @              @       @      @      �?      �?      �?      �?                      �?       @                      @      @      9@       @      @              @       @       @       @                       @      �?      4@      �?       @               @      �?                      (@     �o@     @c@      o@     �a@       @      7@      @      �?      @      �?      @                      �?      @              �?      6@              2@      �?      @              @      �?      �?              �?      �?              n@     �]@      V@      ,@      E@      (@      C@      @     �A@      @      ;@               @      @       @      @              @       @      �?       @                      �?      @              @       @      @                       @      @      @      @      @      �?      @              @      �?      �?      �?                      �?      @                      �?      G@       @      C@               @       @      @       @       @               @       @               @       @              @              c@      Z@      =@      R@      9@      R@       @      @              @       @              1@      Q@      .@      B@      "@     �A@      @      >@      @      4@       @              �?      4@               @      �?      (@              (@      �?                      $@      @      @      @              @      @      @      @      @                      @              �?      @      �?      �?      �?              �?      �?              @               @      @@      �?      @@      �?      ?@      �?      $@              @      �?      @      �?                      @              5@              �?      �?              @              _@      @@      �?       @      �?                       @     �^@      >@     �Q@      @      @      �?      @                      �?      Q@      @      K@      @     �H@       @     �F@      �?      1@              <@      �?      ,@              ,@      �?              �?      ,@              @      �?              �?      @              @       @              �?      @      �?              �?      @              ,@              J@      9@      I@      5@      G@      *@     �@@      *@      $@      "@               @      $@      @              @      $@      @      @      @              �?      @       @       @              �?       @      �?      �?      �?                      �?              �?      @              7@      @      7@      @      $@              *@      @       @              @      @      @                      @              �?      *@              @       @      �?      @      �?      �?      �?                      �?              @      @       @      @                       @       @      @       @      �?              �?       @                      @      @      *@      @      @      @       @      �?       @      �?                       @      @                      @               @r�  tr�  bubhhubehhub.